CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 77 1598 839
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Joe\Documents\School Stuf\Documents\School\Electrical\Circuit Maker 2000 - Portable\BOM.DAT
0 7
2 4 0.500000 0.500000
344 173 457 270
9437202 0
0
6 Title:
5 Name:
0
0
0
332
13 Logic Switch~
5 1118 50 0 10 11
0 564 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3741 0 0
2
41614.3 0
0
13 Logic Switch~
5 1151 46 0 1 11
0 565
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
369 0 0
2
41614.3 1
0
13 Logic Switch~
5 1224 50 0 10 11
0 567 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 S6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8773 0 0
2
41614.3 2
0
13 Logic Switch~
5 1264 51 0 10 11
0 568 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
5 MSBS7
-16 -31 19 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 1 -1 0
1 V
7981 0 0
2
41614.3 3
0
13 Logic Switch~
5 1186 48 0 1 11
0 566
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4205 0 0
2
41614.3 4
0
13 Logic Switch~
5 1084 49 0 1 11
0 563
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 S2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3375 0 0
2
41614.3 5
0
13 Logic Switch~
5 1048 50 0 1 11
0 562
0
0 0 21360 270
2 0V
-6 -21 8 -13
5 LSBS1
-16 -31 19 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
719 0 0
2
41614.3 6
0
9 2-In AND~
219 558 2039 0 3 22
0 6 4 5
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U48D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 23 0
1 U
3749 0 0
2
41614.3 1
0
9 Inverter~
13 628 2062 0 2 22
0 3 6
0
0 0 624 180
6 74LS04
-21 -19 21 -11
5 U128E
-12 -20 23 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 86 0
1 U
3871 0 0
2
41614.3 0
0
9 Inverter~
13 627 1774 0 2 22
0 3 19
0
0 0 624 180
6 74LS04
-21 -19 21 -11
5 U128D
-12 -20 23 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 86 0
1 U
4393 0 0
2
41614.3 0
0
9 2-In AND~
219 557 1751 0 3 22
0 19 12 13
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U48C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 23 0
1 U
6229 0 0
2
41614.3 0
0
8 2-In OR~
219 591 1594 0 3 22
0 3 17 18
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U133B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 91 0
1 U
3757 0 0
2
41614.3 0
0
8 2-In OR~
219 591 1669 0 3 22
0 3 15 16
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U133A
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 91 0
1 U
352 0 0
2
41614.3 0
0
8 2-In OR~
219 594 1867 0 3 22
0 3 11 14
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U132C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 90 0
1 U
3372 0 0
2
41614.3 0
0
8 2-In OR~
219 594 1936 0 3 22
0 3 10 9
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U132B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 90 0
1 U
4911 0 0
2
41614.3 0
0
8 2-In OR~
219 599 2159 0 3 22
0 3 7 8
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U131D
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 89 0
1 U
7574 0 0
2
41614.3 0
0
8 2-In OR~
219 1117 3146 0 3 22
0 3 20 33
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U131C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 89 0
1 U
6601 0 0
2
41614.3 0
0
8 2-In OR~
219 1121 3186 0 3 22
0 596 21 32
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U131B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 89 0
1 U
8531 0 0
2
41614.3 0
0
8 2-In OR~
219 1124 3220 0 3 22
0 3 22 31
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U131A
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 89 0
1 U
6532 0 0
2
41614.3 0
0
8 2-In OR~
219 1126 3260 0 3 22
0 3 23 30
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U130D
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 88 0
1 U
3621 0 0
2
41614.3 0
0
8 2-In OR~
219 1133 3304 0 3 22
0 3 24 29
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U130C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 88 0
1 U
5174 0 0
2
41614.3 0
0
8 2-In OR~
219 1140 3351 0 3 22
0 3 25 28
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U130B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 88 0
1 U
5452 0 0
2
41614.3 0
0
8 2-In OR~
219 1144 3407 0 3 22
0 3 26 27
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U130A
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 88 0
1 U
3626 0 0
2
41614.3 0
0
9 Inverter~
13 3260 3011 0 2 22
0 35 34
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U128C
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 86 0
1 U
3806 0 0
2
5.89641e-315 0
0
5 7415~
219 3271 2954 0 4 22
0 126 127 128 35
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U129A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 87 0
1 U
3389 0 0
2
5.89641e-315 0
0
9 Inverter~
13 3230 3012 0 2 22
0 38 37
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U128B
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 86 0
1 U
9156 0 0
2
5.89641e-315 0
0
9 Inverter~
13 3170 3014 0 2 22
0 39 36
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U128A
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 86 0
1 U
5810 0 0
2
5.89641e-315 0
0
9 Inverter~
13 3086 3012 0 2 22
0 41 40
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126F
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 84 0
1 U
8260 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2995 3010 0 2 22
0 43 42
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126E
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 84 0
1 U
7286 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2906 3010 0 2 22
0 45 44
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126D
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 84 0
1 U
3689 0 0
2
5.89641e-315 0
0
5 7415~
219 3231 2951 0 4 22
0 129 130 131 38
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U127C
16 -3 51 5
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 85 0
1 U
4485 0 0
2
5.89641e-315 0
0
5 7415~
219 3176 2952 0 4 22
0 134 135 136 39
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U127B
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 85 0
1 U
4370 0 0
2
5.89641e-315 0
0
5 7415~
219 3089 2956 0 4 22
0 141 142 143 41
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U127A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 85 0
1 U
7483 0 0
2
5.89641e-315 0
0
5 7415~
219 3001 2956 0 4 22
0 148 149 150 43
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U113A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 67 0
1 U
4214 0 0
2
5.89641e-315 0
0
5 7415~
219 2911 2953 0 4 22
0 48 47 46 45
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U111A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 65 0
1 U
9254 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2820 3005 0 2 22
0 53 52
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126C
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 84 0
1 U
7515 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2726 3004 0 2 22
0 54 49
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126B
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 84 0
1 U
9241 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2650 3000 0 2 22
0 55 50
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U126A
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 84 0
1 U
3783 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2557 2999 0 2 22
0 56 51
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U110A
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 64 0
1 U
5226 0 0
2
5.89641e-315 0
0
5 7415~
219 2817 2952 0 4 22
0 163 164 165 53
0
0 0 624 270
6 74LS15
-21 -28 21 -20
4 U97A
19 -4 47 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 56 0
1 U
6496 0 0
2
5.89641e-315 0
0
5 7415~
219 2732 2954 0 4 22
0 169 170 171 54
0
0 0 624 270
6 74LS15
-21 -28 21 -20
4 U91A
19 -4 47 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 50 0
1 U
6819 0 0
2
5.89641e-315 0
0
5 7415~
219 2652 2952 0 4 22
0 175 176 177 55
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U125C
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 83 0
1 U
6832 0 0
2
5.89641e-315 0
0
5 7415~
219 2561 2947 0 4 22
0 255 256 257 56
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U125B
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 83 0
1 U
7222 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2776 3005 0 2 22
0 58 57
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U123F
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 81 0
1 U
4676 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2687 3006 0 2 22
0 60 59
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U123E
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 81 0
1 U
9334 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2604 3000 0 2 22
0 62 61
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U123D
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 81 0
1 U
4758 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2520 2997 0 2 22
0 64 63
0
0 0 624 270
6 74LS04
-21 -19 21 -11
5 U123C
16 -8 51 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 81 0
1 U
6695 0 0
2
5.89641e-315 0
0
5 7415~
219 2778 2952 0 4 22
0 166 167 168 58
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U125A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 83 0
1 U
8212 0 0
2
5.89641e-315 0
0
5 7415~
219 2694 2951 0 4 22
0 172 173 174 60
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U124C
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 82 0
1 U
3922 0 0
2
5.89641e-315 0
0
5 7415~
219 2609 2948 0 4 22
0 67 66 65 62
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U124B
-3 -7 32 1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 82 0
1 U
7610 0 0
2
5.89641e-315 0
0
5 7415~
219 2522 2945 0 4 22
0 258 259 260 64
0
0 0 624 270
6 74LS15
-21 -28 21 -20
5 U124A
16 -4 51 4
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 82 0
1 U
6131 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2836 259 0 2 22
0 70 71
0
0 0 624 90
6 74LS04
-21 -19 21 -11
5 U123B
16 -2 51 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 81 0
1 U
7187 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2729 257 0 2 22
0 69 72
0
0 0 624 90
6 74LS04
-21 -19 21 -11
5 U123A
16 -2 51 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 81 0
1 U
9198 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2499 265 0 2 22
0 68 73
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U46F
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 22 0
1 U
9468 0 0
2
5.89641e-315 0
0
5 7415~
219 2847 322 0 4 22
0 228 227 226 70
0
0 0 624 90
6 74LS15
-21 -28 21 -20
4 U94A
19 -5 47 3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 53 0
1 U
5160 0 0
2
5.89641e-315 0
0
5 7415~
219 2739 324 0 4 22
0 236 235 234 69
0
0 0 624 90
6 74LS15
-21 -28 21 -20
5 U122C
16 -5 51 3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 3 80 0
1 U
7647 0 0
2
5.89641e-315 0
0
5 7415~
219 2509 332 0 4 22
0 76 75 74 68
0
0 0 624 90
6 74LS15
-21 -28 21 -20
5 U122B
16 -5 51 3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 2 80 0
1 U
7210 0 0
2
5.89641e-315 0
0
9 Inverter~
13 2627 254 0 2 22
0 77 78
0
0 0 624 90
6 74LS04
-21 -19 21 -11
4 U46E
17 -2 45 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 22 0
1 U
7128 0 0
2
5.89641e-315 0
0
5 7415~
219 2637 324 0 4 22
0 243 242 241 77
0
0 0 624 90
6 74LS15
-21 -28 21 -20
5 U122A
16 -5 51 3
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 0 0
65 0 0 0 3 1 80 0
1 U
5367 0 0
2
5.89641e-315 0
0
9 3-In NOR~
219 1698 3241 0 4 22
0 82 88 83 23
0
0 0 624 180
6 74LS27
-21 -24 21 -16
5 U121A
0 -25 35 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 79 0
1 U
7140 0 0
2
5.89641e-315 5.32571e-315
0
9 3-In NOR~
219 1701 3375 0 4 22
0 82 83 84 26
0
0 0 624 180
6 74LS27
-21 -24 21 -16
5 U107C
0 -25 35 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 8 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 3 73 0
1 U
4903 0 0
2
5.89641e-315 5.30499e-315
0
8 4-In OR~
219 1702 3282 0 5 22
0 87 81 86 84 24
0
0 0 624 180
4 4072
-14 -24 14 -16
5 U108B
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 74 0
1 U
3690 0 0
2
5.89641e-315 5.26354e-315
0
9 4-In NOR~
219 1697 3328 0 5 22
0 85 82 86 83 25
0
0 0 624 180
4 4002
-14 -24 14 -16
5 U109B
-4 -25 31 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 2 75 0
1 U
8598 0 0
2
5.89641e-315 0
0
9 Inverter~
13 1696 3204 0 2 22
0 86 22
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U46D
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 22 0
1 U
5737 0 0
2
5.89641e-315 0
0
9 2-In NOR~
219 1696 3169 0 3 22
0 81 89 21
0
0 0 624 180
6 74LS02
-21 -24 21 -16
5 U106D
0 -25 35 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 72 0
1 U
3882 0 0
2
5.89641e-315 0
0
9 2-In NOR~
219 1694 3131 0 3 22
0 88 83 20
0
0 0 624 180
6 74LS02
-21 -24 21 -16
5 U106C
0 -25 35 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 72 0
1 U
3440 0 0
2
5.89641e-315 0
0
8 2-In OR~
219 1946 3447 0 3 22
0 80 99 597
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U120D
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 78 0
1 U
5176 0 0
2
41614.3 7
0
8 2-In OR~
219 1946 3411 0 3 22
0 98 100 87
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U120C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 78 0
1 U
9582 0 0
2
41614.3 8
0
8 2-In OR~
219 1944 3370 0 3 22
0 97 101 82
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U120B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 78 0
1 U
9862 0 0
2
41614.3 9
0
8 2-In OR~
219 1946 3331 0 3 22
0 96 102 81
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U120A
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 78 0
1 U
5432 0 0
2
41614.3 10
0
8 2-In OR~
219 1946 3290 0 3 22
0 95 103 89
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U119D
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 77 0
1 U
3602 0 0
2
41614.3 11
0
8 2-In OR~
219 1946 3249 0 3 22
0 94 104 88
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U119C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 77 0
1 U
4714 0 0
2
41614.3 12
0
8 2-In OR~
219 1947 3210 0 3 22
0 93 105 85
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U119B
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 77 0
1 U
3834 0 0
2
41614.3 13
0
8 2-In OR~
219 1947 3167 0 3 22
0 92 106 86
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U119A
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 77 0
1 U
3577 0 0
2
41614.3 14
0
8 2-In OR~
219 1950 3126 0 3 22
0 91 107 83
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U116D
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 70 0
1 U
7571 0 0
2
41614.3 15
0
8 2-In OR~
219 1948 3088 0 3 22
0 90 108 84
0
0 0 624 180
6 74LS32
-21 -24 21 -16
5 U116C
-6 -25 29 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 70 0
1 U
311 0 0
2
41614.3 16
0
5 7412~
219 3315 2954 0 4 22
0 123 124 125 133
0
0 0 624 270
4 7412
-7 -24 21 -16
5 U118A
17 -7 52 1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 1 76 0
1 U
5524 0 0
2
41614.3 17
0
5 7412~
219 3354 2956 0 4 22
0 120 121 122 132
0
0 0 624 270
4 7412
-7 -24 21 -16
5 U117C
17 -7 52 1
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 6 0
65 0 0 0 3 3 71 0
1 U
6424 0 0
2
41614.3 18
0
8 2-In OR~
219 3333 3011 0 3 22
0 132 133 99
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U116B
26 -7 61 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 70 0
1 U
8878 0 0
2
41614.3 19
0
8 2-In OR~
219 3244 3069 0 3 22
0 34 37 100
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U116A
26 -7 61 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 70 0
1 U
3615 0 0
2
41614.3 20
0
5 7422~
219 3131 2957 0 5 22
0 137 139 138 140 155
0
0 0 624 270
6 74LS22
-21 -28 21 -20
5 U115A
25 -7 60 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 69 0
1 U
7948 0 0
2
41614.3 21
0
8 2-In OR~
219 3154 3065 0 3 22
0 36 155 101
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U112D
28 -7 63 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 66 0
1 U
447 0 0
2
41614.3 22
0
5 7422~
219 3044 2960 0 5 22
0 144 146 145 147 156
0
0 0 624 270
6 74LS22
-21 -28 21 -20
5 U114B
25 -7 60 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 68 0
1 U
4827 0 0
2
41614.3 23
0
8 2-In OR~
219 3065 3059 0 3 22
0 40 156 102
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U112C
28 -7 63 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 66 0
1 U
3675 0 0
2
41614.3 24
0
5 7422~
219 2955 2961 0 5 22
0 151 153 152 154 157
0
0 0 624 270
6 74LS22
-21 -28 21 -20
5 U114A
25 -7 60 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 68 0
1 U
7278 0 0
2
41614.3 25
0
8 2-In OR~
219 2973 3056 0 3 22
0 42 157 103
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U112B
28 -7 63 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 66 0
1 U
926 0 0
2
41614.3 26
0
8 2-In OR~
219 2886 3054 0 3 22
0 44 162 104
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U112A
28 -7 63 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 66 0
1 U
6747 0 0
2
41614.3 27
0
5 7422~
219 2865 2960 0 5 22
0 158 160 159 161 162
0
0 0 624 270
6 74LS22
-21 -28 21 -20
5 U105B
25 -7 60 1
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 63 0
1 U
5177 0 0
2
41614.3 28
0
8 2-In OR~
219 2794 3053 0 3 22
0 52 57 105
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U104D
26 -7 61 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 62 0
1 U
5594 0 0
2
41614.3 29
0
8 2-In OR~
219 2709 3053 0 3 22
0 49 59 106
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U104C
26 -7 61 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 62 0
1 U
9933 0 0
2
41614.3 30
0
8 2-In OR~
219 2625 3050 0 3 22
0 50 61 107
0
0 0 624 270
6 74LS32
-21 -24 21 -16
5 U104B
26 -7 61 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 62 0
1 U
8987 0 0
2
41614.3 31
0
5 7422~
219 3341 318 0 5 22
0 183 181 182 180 209
0
0 0 624 90
6 74LS22
-21 -28 21 -20
5 U105A
23 -2 58 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 63 0
1 U
3275 0 0
2
5.89641e-315 0
0
8 2-In OR~
219 3365 256 0 3 22
0 209 208 80
0
0 0 624 90
6 74LS32
-21 -24 21 -16
5 U104A
26 -3 61 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 62 0
1 U
3551 0 0
2
5.89641e-315 5.26354e-315
0
10 2-In NAND~
219 3389 318 0 3 22
0 179 178 208
0
0 0 624 90
6 74LS00
-14 -24 28 -16
5 U103B
17 -2 52 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 61 0
1 U
9522 0 0
2
5.89641e-315 5.30499e-315
0
5 7422~
219 3250 316 0 5 22
0 189 187 188 186 211
0
0 0 624 90
6 74LS22
-21 -28 21 -20
5 U102B
23 -2 58 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 60 0
1 U
3443 0 0
2
5.89641e-315 5.32571e-315
0
8 2-In OR~
219 3274 254 0 3 22
0 211 210 98
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U99D
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 58 0
1 U
3935 0 0
2
5.89641e-315 5.34643e-315
0
10 2-In NAND~
219 3298 316 0 3 22
0 185 184 210
0
0 0 624 90
6 74LS00
-14 -24 28 -16
5 U103A
17 -2 52 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 61 0
1 U
4532 0 0
2
5.89641e-315 5.3568e-315
0
5 7422~
219 3157 315 0 5 22
0 195 193 194 192 213
0
0 0 624 90
6 74LS22
-21 -28 21 -20
5 U102A
23 -2 58 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 60 0
1 U
7600 0 0
2
5.89641e-315 5.36716e-315
0
8 2-In OR~
219 3181 253 0 3 22
0 213 212 97
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U99C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 58 0
1 U
6952 0 0
2
5.89641e-315 5.37752e-315
0
10 2-In NAND~
219 3205 315 0 3 22
0 191 190 212
0
0 0 624 90
6 74LS00
-14 -24 28 -16
4 U95D
20 -2 48 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 54 0
1 U
3663 0 0
2
5.89641e-315 5.38788e-315
0
5 7422~
219 3064 315 0 5 22
0 201 199 200 198 215
0
0 0 624 90
6 74LS22
-21 -28 21 -20
5 U101B
23 -2 58 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 59 0
1 U
9511 0 0
2
5.89641e-315 5.39306e-315
0
8 2-In OR~
219 3088 253 0 3 22
0 215 214 96
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U99B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 58 0
1 U
4625 0 0
2
5.89641e-315 5.39824e-315
0
10 2-In NAND~
219 3112 315 0 3 22
0 197 196 214
0
0 0 624 90
6 74LS00
-14 -24 28 -16
4 U95C
20 -2 48 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 54 0
1 U
6215 0 0
2
5.89641e-315 5.40342e-315
0
5 7422~
219 2975 317 0 5 22
0 207 205 206 204 217
0
0 0 624 90
6 74LS22
-21 -28 21 -20
5 U101A
23 -2 58 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 59 0
1 U
4535 0 0
2
5.89641e-315 5.4086e-315
0
8 2-In OR~
219 2999 255 0 3 22
0 217 216 95
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U99A
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 58 0
1 U
3611 0 0
2
5.89641e-315 5.41378e-315
0
10 2-In NAND~
219 3023 317 0 3 22
0 203 202 216
0
0 0 624 90
6 74LS00
-14 -24 28 -16
4 U95B
20 -2 48 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 54 0
1 U
9183 0 0
2
5.89641e-315 5.41896e-315
0
10 2-In NAND~
219 2933 319 0 3 22
0 219 218 224
0
0 0 624 90
6 74LS00
-14 -24 28 -16
4 U95A
20 -2 48 6
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 54 0
1 U
3593 0 0
2
5.89641e-315 5.42414e-315
0
8 2-In OR~
219 2909 257 0 3 22
0 225 224 94
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U96D
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 55 0
1 U
4142 0 0
2
5.89641e-315 5.42933e-315
0
5 7422~
219 2885 319 0 5 22
0 223 221 222 220 225
0
0 0 624 90
6 74LS22
-21 -28 21 -20
4 U98B
26 -2 54 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 57 0
1 U
9564 0 0
2
5.89641e-315 5.43192e-315
0
5 7422~
219 2796 320 0 5 22
0 232 230 231 229 233
0
0 0 624 90
6 74LS22
-21 -28 21 -20
4 U98A
26 -2 54 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 57 0
1 U
7772 0 0
2
5.89641e-315 5.4371e-315
0
8 2-In OR~
219 2815 194 0 3 22
0 233 71 93
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U96C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 55 0
1 U
3826 0 0
2
5.89641e-315 5.43969e-315
0
5 7422~
219 2688 321 0 5 22
0 240 238 239 237 248
0
0 0 624 90
6 74LS22
-21 -28 21 -20
4 U93B
26 -2 54 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 52 0
1 U
9216 0 0
2
5.89641e-315 5.44487e-315
0
8 2-In OR~
219 2714 196 0 3 22
0 248 72 92
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U92D
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 51 0
1 U
770 0 0
2
5.89641e-315 5.44746e-315
0
5 7422~
219 2585 321 0 5 22
0 247 245 246 244 249
0
0 0 624 90
6 74LS22
-21 -28 21 -20
4 U93A
26 -2 54 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 52 0
1 U
6894 0 0
2
5.89641e-315 5.45264e-315
0
8 2-In OR~
219 2608 196 0 3 22
0 249 78 91
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U92C
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 51 0
1 U
3840 0 0
2
5.89641e-315 5.45523e-315
0
8 2-In OR~
219 2482 198 0 3 22
0 250 73 90
0
0 0 624 90
6 74LS32
-21 -24 21 -16
4 U92B
29 -3 57 5
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 51 0
1 U
6568 0 0
2
5.89641e-315 5.45782e-315
0
5 7422~
219 2458 327 0 5 22
0 254 252 253 251 250
0
0 0 624 90
6 74LS22
-21 -28 21 -20
4 U89A
26 -2 54 6
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 48 0
1 U
656 0 0
2
5.89641e-315 5.46041e-315
0
7 74LS154
95 2941 1069 0 22 45
0 116 116 119 79 118 117 206 222 231
239 246 253 183 189 195 201 207 223 232
240 247 254
0
0 0 4848 602
7 74LS154
-24 -87 25 -79
4 U100
84 -3 112 5
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
5430 0 0
2
5.89641e-315 5.46559e-315
0
7 74LS154
95 3091 1069 0 22 45
0 115 115 119 79 118 117 244 251 181
187 193 199 205 221 230 238 245 252 182
188 194 200
0
0 0 4848 602
7 74LS154
-24 -87 25 -79
3 U90
83 -3 104 5
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
6853 0 0
2
5.89641e-315 5.46818e-315
0
7 74LS154
95 3237 1069 0 22 45
0 114 114 119 79 118 117 191 197 203
219 228 236 243 76 180 186 192 198 204
220 229 237
0
0 0 4848 602
7 74LS154
-24 -87 25 -79
3 U87
83 -3 104 5
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3322 0 0
2
5.89641e-315 5.47077e-315
0
7 74LS154
95 3384 1070 0 22 45
0 113 113 119 79 118 117 226 234 241
74 178 184 190 196 202 218 227 235 242
75 179 185
0
0 0 4848 602
7 74LS154
-24 -87 25 -79
3 U88
83 -3 104 5
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
9236 0 0
2
5.89641e-315 5.47207e-315
0
8 2-In OR~
219 2537 3045 0 3 22
0 51 63 108
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U92A
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 51 0
1 U
8728 0 0
2
5.89641e-315 5.47336e-315
0
7 74LS154
95 3240 2196 0 22 45
0 110 110 119 79 118 117 176 256 121
127 136 143 150 46 165 171 177 257 122
128 137 144
0
0 0 4848 270
7 74LS154
-24 -87 25 -79
3 U86
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
4790 0 0
2
5.89641e-315 5.47725e-315
0
7 74LS154
95 3387 2197 0 22 45
0 109 109 119 79 118 117 134 141 148
48 163 169 175 255 120 126 135 142 149
47 164 170
0
0 0 4848 270
7 74LS154
-24 -87 25 -79
3 U85
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3447 0 0
2
5.89641e-315 5.47854e-315
0
7 74LS154
95 3094 2196 0 22 45
0 111 111 119 79 118 117 151 158 166
172 67 258 123 129 138 145 152 159 167
173 66 259
0
0 0 4848 270
7 74LS154
-24 -87 25 -79
3 U84
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
4769 0 0
2
5.89641e-315 5.47984e-315
0
7 74LS154
95 2944 2196 0 22 45
0 112 112 119 79 118 117 124 130 139
146 153 160 168 174 65 260 125 131 140
147 154 161
0
0 0 4848 270
7 74LS154
-24 -87 25 -79
3 U82
83 -2 104 6
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3989 0 0
2
5.89641e-315 5.48113e-315
0
9 4-In NOR~
219 898 2009 0 5 22
0 263 264 265 262 4
0
0 0 624 180
4 4002
-14 -24 14 -16
5 U109A
-4 -25 31 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
11 typeDigital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 9 0
65 0 0 0 2 1 75 0
1 U
3188 0 0
2
41614.3 32
0
8 4-In OR~
219 900 1907 0 5 22
0 266 267 265 261 10
0
0 0 624 180
4 4072
-14 -24 14 -16
5 U108A
-10 -25 25 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 74 0
1 U
7596 0 0
2
41614.3 33
0
9 3-In NOR~
219 900 2122 0 4 22
0 263 262 261 7
0
0 0 624 180
6 74LS27
-21 -24 21 -16
5 U107B
0 -25 35 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 2 73 0
1 U
4823 0 0
2
41614.3 34
0
9 3-In NOR~
219 896 1841 0 4 22
0 263 268 262 11
0
0 0 624 180
6 74LS27
-21 -24 21 -16
5 U107A
0 -25 35 -17
0
15 DVCC=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 13 12 1 2 13 12 3
4 5 6 9 10 11 8 0 0 0
0 6 0
65 0 0 0 3 1 73 0
1 U
8750 0 0
2
41614.3 35
0
9 Inverter~
13 892 1718 0 2 22
0 265 12
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U46C
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 22 0
1 U
8804 0 0
2
41614.3 36
0
9 2-In NOR~
219 894 1646 0 3 22
0 267 269 15
0
0 0 624 180
6 74LS02
-21 -24 21 -16
5 U106B
0 -25 35 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 72 0
1 U
9238 0 0
2
41614.3 37
0
9 2-In NOR~
219 898 1571 0 3 22
0 268 262 17
0
0 0 624 180
6 74LS02
-21 -24 21 -16
5 U106A
0 -25 35 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 72 0
1 U
8829 0 0
2
41614.3 38
0
8 2-In OR~
219 1154 1789 0 3 22
0 272 274 265
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U81D
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 47 0
1 U
4267 0 0
2
41614.3 39
0
8 2-In OR~
219 1149 1663 0 3 22
0 271 275 262
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U81C
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 47 0
1 U
4134 0 0
2
41614.3 40
0
8 2-In OR~
219 1151 1539 0 3 22
0 270 276 261
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U81B
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 47 0
1 U
9687 0 0
2
41614.3 41
0
8 2-In OR~
219 1245 3015 0 3 22
0 273 278 272
0
0 0 624 180
6 74LS32
-21 -24 21 -16
4 U81A
-2 -25 26 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 47 0
1 U
3640 0 0
2
5.89641e-315 5.48243e-315
0
5 7422~
219 1355 2971 0 5 22
0 283 285 284 286 278
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U83B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 49 0
1 U
3203 0 0
2
5.89641e-315 5.48372e-315
0
5 7422~
219 1356 3018 0 5 22
0 279 281 280 282 273
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U83A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 49 0
1 U
3606 0 0
2
5.89641e-315 5.48502e-315
0
5 7422~
219 1349 2846 0 5 22
0 293 295 294 296 409
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U80B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 46 0
1 U
6649 0 0
2
5.89641e-315 5.48631e-315
0
5 7422~
219 1350 2893 0 5 22
0 289 291 290 292 408
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U80A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 46 0
1 U
3797 0 0
2
5.89641e-315 5.48761e-315
0
10 2-In NAND~
219 1352 2932 0 3 22
0 287 288 407
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U75D
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 41 0
1 U
7609 0 0
2
5.89641e-315 5.4889e-315
0
8 3-In OR~
219 1247 2891 0 4 22
0 407 408 409 271
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U77C
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 43 0
1 U
5110 0 0
2
5.89641e-315 5.4902e-315
0
5 7422~
219 1346 2722 0 5 22
0 303 305 304 306 412
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U79B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 45 0
1 U
9643 0 0
2
5.89641e-315 5.49149e-315
0
5 7422~
219 1347 2769 0 5 22
0 299 301 300 302 411
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U79A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 45 0
1 U
3480 0 0
2
5.89641e-315 5.49279e-315
0
10 2-In NAND~
219 1349 2808 0 3 22
0 297 298 410
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U75C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 41 0
1 U
3609 0 0
2
5.89641e-315 5.49408e-315
0
8 3-In OR~
219 1244 2767 0 4 22
0 410 411 412 270
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U77B
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 43 0
1 U
8185 0 0
2
5.89641e-315 5.49538e-315
0
5 7422~
219 1346 2597 0 5 22
0 313 315 314 316 415
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U78B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 44 0
1 U
5744 0 0
2
5.89641e-315 5.49667e-315
0
5 7422~
219 1347 2644 0 5 22
0 309 311 310 312 414
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U78A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 44 0
1 U
9374 0 0
2
5.89641e-315 5.49797e-315
0
10 2-In NAND~
219 1349 2683 0 3 22
0 307 308 413
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U75B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 41 0
1 U
7786 0 0
2
5.89641e-315 5.49926e-315
0
8 3-In OR~
219 1244 2642 0 4 22
0 413 414 415 598
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U77A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 512 3 1 43 0
1 U
6749 0 0
2
5.89641e-315 5.50056e-315
0
5 7422~
219 1344 2471 0 5 22
0 323 325 324 326 418
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U76B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 42 0
1 U
4813 0 0
2
5.89641e-315 5.50185e-315
0
5 7422~
219 1345 2518 0 5 22
0 319 321 320 322 417
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U76A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 42 0
1 U
4826 0 0
2
5.89641e-315 5.50315e-315
0
10 2-In NAND~
219 1347 2557 0 3 22
0 317 318 416
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U75A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 41 0
1 U
765 0 0
2
5.89641e-315 5.50444e-315
0
8 3-In OR~
219 1242 2516 0 4 22
0 416 417 418 266
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U72C
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 38 0
1 U
6493 0 0
2
5.89641e-315 5.50574e-315
0
5 7422~
219 1339 2346 0 5 22
0 333 335 334 336 421
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U74B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 40 0
1 U
9234 0 0
2
5.89641e-315 5.50703e-315
0
5 7422~
219 1340 2393 0 5 22
0 329 331 330 332 420
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U74A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 40 0
1 U
8902 0 0
2
5.89641e-315 5.50833e-315
0
10 2-In NAND~
219 1342 2432 0 3 22
0 327 328 419
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U69D
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 35 0
1 U
596 0 0
2
5.89641e-315 5.50963e-315
0
8 3-In OR~
219 1237 2391 0 4 22
0 419 420 421 263
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U72B
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 38 0
1 U
5799 0 0
2
5.89641e-315 5.51092e-315
0
5 7422~
219 1336 2225 0 5 22
0 343 345 344 346 424
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U73B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 39 0
1 U
4948 0 0
2
5.89641e-315 5.51222e-315
0
5 7422~
219 1337 2272 0 5 22
0 339 341 340 342 423
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U73A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 39 0
1 U
3151 0 0
2
5.89641e-315 5.51286e-315
0
10 2-In NAND~
219 1339 2311 0 3 22
0 337 338 422
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U69C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 35 0
1 U
7543 0 0
2
5.89641e-315 5.51351e-315
0
8 3-In OR~
219 1234 2270 0 4 22
0 422 423 424 267
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U72A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 38 0
1 U
3946 0 0
2
5.89641e-315 5.51416e-315
0
5 7422~
219 1332 2098 0 5 22
0 353 355 354 356 427
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U71B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 37 0
1 U
8784 0 0
2
5.89641e-315 5.51481e-315
0
5 7422~
219 1333 2145 0 5 22
0 349 351 350 352 426
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U71A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 37 0
1 U
3459 0 0
2
5.89641e-315 5.51545e-315
0
10 2-In NAND~
219 1335 2184 0 3 22
0 347 348 425
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U69B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 35 0
1 U
9264 0 0
2
5.89641e-315 5.5161e-315
0
8 3-In OR~
219 1230 2143 0 4 22
0 425 426 427 269
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U67C
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 33 0
1 U
422 0 0
2
5.89641e-315 5.51675e-315
0
5 7422~
219 1328 1976 0 5 22
0 363 365 364 366 430
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U70B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 36 0
1 U
5301 0 0
2
5.89641e-315 5.5174e-315
0
5 7422~
219 1329 2023 0 5 22
0 359 361 360 362 429
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U70A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 36 0
1 U
3416 0 0
2
5.89641e-315 5.51804e-315
0
10 2-In NAND~
219 1331 2062 0 3 22
0 357 358 428
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U69A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 35 0
1 U
8994 0 0
2
5.89641e-315 5.51869e-315
0
8 3-In OR~
219 1226 2021 0 4 22
0 428 429 430 268
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U67B
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 33 0
1 U
4927 0 0
2
5.89641e-315 5.51934e-315
0
5 7422~
219 1324 1851 0 5 22
0 373 375 374 376 433
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U68B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 34 0
1 U
3312 0 0
2
5.89641e-315 5.51999e-315
0
5 7422~
219 1325 1898 0 5 22
0 369 371 370 372 432
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U68A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 34 0
1 U
8964 0 0
2
5.89641e-315 5.52063e-315
0
10 2-In NAND~
219 1327 1937 0 3 22
0 367 368 431
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U63D
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 29 0
1 U
4138 0 0
2
5.89641e-315 5.52128e-315
0
8 3-In OR~
219 1222 1896 0 4 22
0 431 432 433 264
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U67A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 33 0
1 U
392 0 0
2
5.89641e-315 5.52193e-315
0
5 7422~
219 1321 1731 0 5 22
0 383 385 384 386 436
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U66B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 32 0
1 U
4526 0 0
2
5.89641e-315 5.52258e-315
0
5 7422~
219 1322 1778 0 5 22
0 379 381 380 382 435
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U66A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 32 0
1 U
6971 0 0
2
5.89641e-315 5.52322e-315
0
10 2-In NAND~
219 1324 1817 0 3 22
0 377 378 434
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U63C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
4845 0 0
2
5.89641e-315 5.52387e-315
0
8 3-In OR~
219 1219 1776 0 4 22
0 434 435 436 274
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U64C
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 30 0
1 U
7679 0 0
2
5.89641e-315 5.52452e-315
0
5 7422~
219 1320 1605 0 5 22
0 393 395 394 396 439
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U65B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 31 0
1 U
3883 0 0
2
5.89641e-315 5.52517e-315
0
5 7422~
219 1321 1652 0 5 22
0 389 391 390 392 438
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U65A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 31 0
1 U
3876 0 0
2
5.89641e-315 5.52581e-315
0
10 2-In NAND~
219 1323 1691 0 3 22
0 387 388 437
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U63B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 29 0
1 U
6399 0 0
2
5.89641e-315 5.52646e-315
0
8 3-In OR~
219 1218 1650 0 4 22
0 437 438 439 275
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U64B
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 30 0
1 U
3299 0 0
2
5.89641e-315 5.52711e-315
0
8 3-In OR~
219 1215 1520 0 4 22
0 440 441 442 276
0
0 0 624 180
4 4075
-14 -24 14 -16
4 U64A
-2 -25 26 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 30 0
1 U
8181 0 0
2
5.89641e-315 5.52776e-315
0
10 2-In NAND~
219 1320 1561 0 3 22
0 397 398 440
0
0 0 624 180
6 74LS00
-14 -24 28 -16
4 U63A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
3458 0 0
2
5.89641e-315 5.52841e-315
0
5 7422~
219 1318 1522 0 5 22
0 399 401 400 402 441
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U62B
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 13 12 10 9 8 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 2 28 0
1 U
899 0 0
2
5.89641e-315 5.52905e-315
0
5 7422~
219 1317 1475 0 5 22
0 403 405 404 406 442
0
0 0 624 180
6 74LS22
-21 -28 21 -20
4 U62A
-11 -31 17 -23
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 13 12 10 9 8 0 0 0 0
0 0 0
65 0 0 0 2 1 28 0
1 U
4812 0 0
2
5.89641e-315 5.5297e-315
0
8 4-In OR~
219 1766 2753 0 5 22
0 443 444 453 3 109
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U61A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 27 0
1 U
3617 0 0
2
41614.3 42
0
8 4-In OR~
219 1762 2593 0 5 22
0 446 444 453 3 110
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U60B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 26 0
1 U
9290 0 0
2
41614.3 43
0
8 4-In OR~
219 1758 2424 0 5 22
0 443 447 453 3 111
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U60A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 26 0
1 U
5248 0 0
2
41614.3 44
0
8 4-In OR~
219 1756 2266 0 5 22
0 446 447 453 3 112
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U59B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 25 0
1 U
8646 0 0
2
41614.3 45
0
8 4-In OR~
219 1753 2096 0 5 22
0 443 444 445 3 113
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U59A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 25 0
1 U
6620 0 0
2
41614.3 46
0
8 4-In OR~
219 1751 1933 0 5 22
0 446 444 445 3 114
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U58B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 24 0
1 U
6104 0 0
2
41614.3 47
0
8 4-In OR~
219 1748 1772 0 5 22
0 443 447 445 3 115
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U58A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 24 0
1 U
3235 0 0
2
41614.3 48
0
8 4-In OR~
219 1746 1608 0 5 22
0 446 447 445 3 116
0
0 0 624 180
4 4072
-14 -24 14 -16
4 U31B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 19 0
1 U
4598 0 0
2
41614.3 49
0
7 74LS154
95 1615 2195 0 22 45
0 112 112 119 79 118 117 327 328 329
330 331 332 333 334 335 336 337 338 339
340 341 342
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U57
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
4385 0 0
2
41614.3 50
0
7 74LS154
95 1616 2358 0 22 45
0 111 111 119 79 118 117 311 312 313
314 315 316 317 318 319 320 321 322 323
324 325 326
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U56
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
8444 0 0
2
41614.3 51
0
7 74LS154
95 1617 2686 0 22 45
0 109 109 119 79 118 117 279 280 281
282 283 284 285 286 287 288 289 290 291
292 293 294
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U55
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3718 0 0
2
41614.3 52
0
7 74LS154
95 1616 2523 0 22 45
0 110 110 119 79 118 117 295 296 297
298 299 300 301 302 303 304 305 306 307
308 309 310
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U54
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
9950 0 0
2
41614.3 53
0
7 74LS154
95 1615 1864 0 22 45
0 114 114 119 79 118 117 359 360 361
362 363 364 365 366 367 368 369 370 371
372 373 374
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U53
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
4505 0 0
2
41614.3 54
0
7 74LS154
95 1616 2027 0 22 45
0 113 113 119 79 118 117 343 344 345
346 347 348 349 350 351 352 353 354 355
356 357 358
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U52
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3627 0 0
2
41614.3 55
0
7 74LS154
95 1615 1699 0 22 45
0 115 115 119 79 118 117 375 376 377
378 379 380 381 382 383 384 385 386 387
388 389 390
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U51
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
3310 0 0
2
41614.3 56
0
7 74LS154
95 1614 1536 0 22 45
0 116 116 119 79 118 117 391 392 393
394 395 396 397 398 399 400 401 402 403
404 405 406
0
0 0 4848 180
7 74LS154
-24 -87 25 -79
3 U50
-11 -88 10 -80
0
16 DVCC=24;DGND=12;
155 %D [%24bi %12bi %1i %2i %3i %4i %5i %6i]
+ [%24bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o %19o %20o %21o %22o] %M
0
12 type:digital
5 DIP24
45

0 19 18 20 21 22 23 17 16 15
14 13 11 10 9 8 7 6 5 4
3 2 1 19 18 20 21 22 23 17
16 15 14 13 11 10 9 8 7 6
5 4 3 2 1 0
65 0 0 0 1 0 0 0
1 U
474 0 0
2
41614.3 57
0
13 SR Flip-Flop~
219 2856 917 0 4 9
0 463 462 454 3
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U49
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7310 0 0
2
5.89641e-315 5.53035e-315
0
9 2-In AND~
219 2821 817 0 3 22
0 452 464 462
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U48B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 23 0
1 U
9609 0 0
2
5.89641e-315 5.531e-315
0
9 2-In AND~
219 2884 818 0 3 22
0 448 452 463
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U48A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 23 0
1 U
7364 0 0
2
5.89641e-315 5.53164e-315
0
9 Inverter~
13 2809 739 0 2 22
0 448 464
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U46B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 22 0
1 U
3943 0 0
2
5.89641e-315 5.53229e-315
0
13 SR Flip-Flop~
219 2742 915 0 4 9
0 466 465 453 445
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U47
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3496 0 0
2
5.89641e-315 5.53294e-315
0
9 2-In AND~
219 2707 815 0 3 22
0 452 467 465
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U44D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 21 0
1 U
7335 0 0
2
5.89641e-315 5.53359e-315
0
9 2-In AND~
219 2770 816 0 3 22
0 449 452 466
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U44C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 21 0
1 U
458 0 0
2
5.89641e-315 5.53423e-315
0
9 Inverter~
13 2695 737 0 2 22
0 449 467
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U46A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 22 0
1 U
6142 0 0
2
5.89641e-315 5.53488e-315
0
13 SR Flip-Flop~
219 2625 917 0 4 9
0 469 468 444 447
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U45
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9664 0 0
2
5.89641e-315 5.53553e-315
0
9 2-In AND~
219 2590 817 0 3 22
0 452 470 468
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U44B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 21 0
1 U
9203 0 0
2
5.89641e-315 5.53618e-315
0
9 2-In AND~
219 2653 818 0 3 22
0 450 452 469
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U44A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 21 0
1 U
3372 0 0
2
5.89641e-315 5.53682e-315
0
9 Inverter~
13 2578 739 0 2 22
0 450 470
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 16 0
1 U
5771 0 0
2
5.89641e-315 5.53747e-315
0
13 SR Flip-Flop~
219 2508 918 0 4 9
0 472 471 443 446
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U43
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
3554 0 0
2
5.89641e-315 5.53812e-315
0
9 2-In AND~
219 2473 818 0 3 22
0 452 473 471
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U41D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 20 0
1 U
3823 0 0
2
5.89641e-315 5.53877e-315
0
9 2-In AND~
219 2536 819 0 3 22
0 451 452 472
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U41C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 20 0
1 U
6185 0 0
2
5.89641e-315 5.53941e-315
0
9 Inverter~
13 2461 740 0 2 22
0 451 473
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 16 0
1 U
4465 0 0
2
5.89641e-315 5.54006e-315
0
13 SR Flip-Flop~
219 2401 919 0 4 9
0 475 474 457 119
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U42
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
9574 0 0
2
5.89641e-315 5.54071e-315
0
9 2-In AND~
219 2366 819 0 3 22
0 452 476 474
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U41B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 20 0
1 U
7277 0 0
2
5.89641e-315 5.54136e-315
0
9 2-In AND~
219 2429 820 0 3 22
0 277 452 475
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U41A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 20 0
1 U
7450 0 0
2
5.89641e-315 5.542e-315
0
9 Inverter~
13 2354 741 0 2 22
0 277 476
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 16 0
1 U
3892 0 0
2
5.89641e-315 5.54265e-315
0
13 SR Flip-Flop~
219 2291 917 0 4 9
0 478 477 455 79
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U40
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
5444 0 0
2
5.89641e-315 5.5433e-315
0
9 2-In AND~
219 2256 817 0 3 22
0 452 479 477
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U38D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 17 0
1 U
777 0 0
2
5.89641e-315 5.54395e-315
0
9 2-In AND~
219 2319 818 0 3 22
0 459 452 478
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U38C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 17 0
1 U
3280 0 0
2
5.89641e-315 5.54459e-315
0
9 Inverter~
13 2244 739 0 2 22
0 459 479
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 16 0
1 U
5774 0 0
2
5.89641e-315 5.54524e-315
0
13 SR Flip-Flop~
219 2183 915 0 4 9
0 481 480 456 118
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U39
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
5917 0 0
2
5.89641e-315 5.54589e-315
0
9 2-In AND~
219 2148 815 0 3 22
0 452 482 480
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U38B
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 17 0
1 U
5823 0 0
2
5.89641e-315 5.54654e-315
0
9 2-In AND~
219 2211 816 0 3 22
0 460 452 481
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U38A
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 17 0
1 U
3536 0 0
2
5.89641e-315 5.54719e-315
0
9 Inverter~
13 2136 737 0 2 22
0 460 482
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 16 0
1 U
3383 0 0
2
5.89641e-315 5.54783e-315
0
9 Inverter~
13 2016 739 0 2 22
0 461 485
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U37A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 16 0
1 U
331 0 0
2
5.89641e-315 5.54848e-315
0
9 2-In AND~
219 2091 818 0 3 22
0 461 452 484
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U35D
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 15 0
1 U
9968 0 0
2
5.89641e-315 5.54913e-315
0
9 2-In AND~
219 2028 817 0 3 22
0 452 485 483
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U35C
17 -4 45 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
7505 0 0
2
5.89641e-315 5.54978e-315
0
13 SR Flip-Flop~
219 2063 917 0 4 9
0 484 483 458 117
0
0 0 4720 270
4 SRFF
-14 -53 14 -45
3 U36
24 -34 45 -26
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
7962 0 0
2
5.89641e-315 5.55042e-315
0
9 Inverter~
13 1968 133 0 2 22
0 489 490
0
0 0 624 180
6 74LS04
-21 -19 21 -11
4 U24F
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 11 0
1 U
3622 0 0
2
5.89641e-315 5.55107e-315
0
9 2-In AND~
219 1900 165 0 3 22
0 489 452 488
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U35B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
4473 0 0
2
5.89641e-315 5.55172e-315
0
9 2-In AND~
219 1902 127 0 3 22
0 490 452 487
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U35A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
4493 0 0
2
5.89641e-315 5.55237e-315
0
13 SR Flip-Flop~
219 1815 182 0 4 9
0 488 487 599 486
0
0 0 4720 512
4 SRFF
-14 -53 14 -45
3 U32
-6 -55 15 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
6230 0 0
2
5.89641e-315 5.55301e-315
0
4 4585
219 2111 382 0 14 29
0 2 491 491 2 448 449 450 451 494
493 492 600 601 489
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U34
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
6181 0 0
2
41614.3 58
0
4 4585
219 2022 261 0 14 29
0 2 491 2 2 277 459 460 461 602
491 603 492 493 494
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U30
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
3165 0 0
2
41614.3 59
0
14 Logic Display~
6 769 211 0 1 2
46 452
0
0 0 53856 0
6 100MEG
3 -16 45 -8
4 STOP
-15 -21 13 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7499 0 0
2
41614.3 60
0
14 Logic Display~
6 743 213 0 1 2
45 496
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 GO
-8 -23 6 -15
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8986 0 0
2
41614.3 61
0
9 CC 7-Seg~
183 662 209 0 17 19
10 33 32 31 30 29 28 27 604 2
1 1 1 1 1 1 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP3
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3568 0 0
2
41614.3 62
0
9 CC 7-Seg~
183 602 211 0 17 19
10 18 16 13 14 9 5 8 605 2
1 1 1 1 1 1 0 2
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
8397 0 0
2
41614.3 63
0
9 CC 7-Seg~
183 541 212 0 17 19
10 486 491 491 486 486 486 2 491 2
1 1 1 1 1 1 0 1
0
0 0 20576 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 0 1 0 0 0
4 DISP
311 0 0
2
41614.3 64
0
7 Buffer~
58 543 15 0 2 22
0 497 498
0
0 0 624 0
4 4050
-14 -19 14 -11
4 U27F
-14 -20 14 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 12 0
1 U
3832 0 0
2
41614.3 65
0
9 2-In AND~
219 1042 1129 0 3 22
0 497 510 506
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U29D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3263 0 0
2
5.89641e-315 5.55366e-315
0
9 2-In AND~
219 1045 1427 0 3 22
0 497 507 499
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U29C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
4814 0 0
2
5.89641e-315 5.55398e-315
0
9 2-In AND~
219 1040 1380 0 3 22
0 497 519 500
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U29B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
3278 0 0
2
5.89641e-315 5.55431e-315
0
9 2-In AND~
219 1040 1336 0 3 22
0 497 508 501
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U29A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6768 0 0
2
5.89641e-315 5.55463e-315
0
9 2-In AND~
219 1040 1293 0 3 22
0 497 520 502
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U28D
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 13 0
1 U
3687 0 0
2
5.89641e-315 5.55496e-315
0
9 2-In AND~
219 1040 1251 0 3 22
0 497 521 503
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U28C
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 13 0
1 U
4404 0 0
2
5.89641e-315 5.55528e-315
0
9 2-In AND~
219 1040 1212 0 3 22
0 497 509 504
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U28B
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 13 0
1 U
3705 0 0
2
5.89641e-315 5.5556e-315
0
9 2-In AND~
219 1040 1170 0 3 22
0 522 497 505
0
0 0 624 180
6 74LS08
-21 -24 21 -16
4 U28A
-16 -25 12 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 13 0
1 U
5509 0 0
2
5.89641e-315 5.55593e-315
0
7 Buffer~
58 778 731 0 2 22
0 512 511
0
0 0 624 0
4 4050
-14 -19 14 -11
4 U27E
-14 -20 14 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 5 12 0
1 U
6447 0 0
2
5.89641e-315 5.55625e-315
0
7 Buffer~
58 603 710 0 2 22
0 514 513
0
0 0 624 0
4 4050
-14 -19 14 -11
4 U27D
-14 -20 14 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 12 0
1 U
3260 0 0
2
5.89641e-315 5.55657e-315
0
7 Buffer~
58 643 450 0 2 22
0 499 515
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U27C
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 12 0
1 U
7932 0 0
2
5.89641e-315 5.5569e-315
0
7 Buffer~
58 580 447 0 2 22
0 500 517
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U27B
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 12 0
1 U
3293 0 0
2
5.89641e-315 5.55722e-315
0
9 Inverter~
13 593 529 0 2 22
0 517 518
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U24E
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 11 0
1 U
4463 0 0
2
5.89641e-315 5.55755e-315
0
9 2-In AND~
219 578 583 0 3 22
0 518 517 514
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11D
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 7 0
1 U
3841 0 0
2
5.89641e-315 5.55787e-315
0
9 Inverter~
13 656 531 0 2 22
0 515 516
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U24D
13 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 11 0
1 U
7621 0 0
2
5.89641e-315 5.55819e-315
0
9 2-In AND~
219 641 585 0 3 22
0 516 515 512
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11C
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 7 0
1 U
3390 0 0
2
5.89641e-315 5.55852e-315
0
7 Buffer~
58 1542 977 0 2 22
0 523 510
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U27A
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 12 0
1 U
96 0 0
2
5.89641e-315 5.55884e-315
0
7 Buffer~
58 1515 976 0 2 22
0 524 522
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U22F
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 10 0
1 U
3532 0 0
2
5.89641e-315 5.55917e-315
0
7 Buffer~
58 1489 978 0 2 22
0 525 509
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U22E
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 5 10 0
1 U
3134 0 0
2
5.89641e-315 5.55949e-315
0
7 Buffer~
58 1465 977 0 2 22
0 526 521
0
0 0 624 270
4 4050
-14 -19 14 -11
4 U22D
14 -5 42 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 10 0
1 U
5510 0 0
2
5.89641e-315 5.55981e-315
0
6 74LS83
105 1633 959 0 14 29
0 2 2 2 2 530 529 528 527 531
507 519 508 520 606
0
0 0 4848 782
6 74LS83
-21 -60 21 -52
3 U26
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3430 0 0
2
5.89641e-315 5.56014e-315
0
6 74LS83
105 1507 829 0 14 29
0 2 2 2 2 535 534 533 532 491
526 525 524 523 531
0
0 0 4848 782
6 74LS83
-21 -60 21 -52
3 U25
56 -2 77 6
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
999 0 0
2
5.89641e-315 5.56046e-315
0
9 Inverter~
13 1629 679 0 2 22
0 451 527
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U24C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 11 0
1 U
6527 0 0
2
5.89641e-315 5.56078e-315
0
9 Inverter~
13 1668 678 0 2 22
0 450 528
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U24B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 11 0
1 U
6717 0 0
2
5.89641e-315 5.56111e-315
0
9 Inverter~
13 1705 674 0 2 22
0 449 529
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U24A
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
5410 0 0
2
5.89641e-315 5.56143e-315
0
9 Inverter~
13 1745 676 0 2 22
0 448 530
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U20F
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 9 0
1 U
8250 0 0
2
5.89641e-315 5.56176e-315
0
9 Inverter~
13 1544 674 0 2 22
0 459 534
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U20E
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 9 0
1 U
327 0 0
2
5.89641e-315 5.56208e-315
0
9 Inverter~
13 1584 676 0 2 22
0 277 535
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U20D
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 9 0
1 U
3833 0 0
2
5.89641e-315 5.5624e-315
0
9 Inverter~
13 1507 678 0 2 22
0 460 533
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U20C
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 9 0
1 U
3474 0 0
2
5.89641e-315 5.56273e-315
0
9 Inverter~
13 1467 676 0 2 22
0 461 532
0
0 0 624 270
6 74LS04
-21 -19 21 -11
4 U20B
17 -8 45 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 9 0
1 U
9900 0 0
2
5.89641e-315 5.56305e-315
0
8 4-In OR~
219 186 190 0 5 22
0 506 536 538 539 540
0
0 0 624 270
4 4072
-14 -24 14 -16
4 U31A
27 -5 55 3
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 19 0
1 U
9419 0 0
2
41614.3 66
0
8 3-In OR~
219 388 183 0 4 22
0 503 536 541 542
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U33C
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 18 0
1 U
6151 0 0
2
41614.3 67
0
8 3-In OR~
219 246 166 0 4 22
0 505 537 541 543
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U33B
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 18 0
1 U
3237 0 0
2
41614.3 68
0
8 2-In OR~
219 314 163 0 3 22
0 504 538 544
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U12D
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 8 0
1 U
7123 0 0
2
41614.3 69
0
8 2-In OR~
219 494 433 0 3 22
0 501 537 580
0
0 0 624 270
6 74LS32
-21 -24 21 -16
4 U12C
29 -7 57 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 8 0
1 U
4133 0 0
2
41614.3 70
0
8 3-In OR~
219 431 433 0 4 22
0 502 537 536 545
0
0 0 624 270
4 4075
-14 -24 14 -16
4 U33A
29 -7 57 1
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 18 0
1 U
3640 0 0
2
41614.3 71
0
12 D Flip-Flop~
219 1251 663 0 4 9
0 547 546 607 448
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U23
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
9534 0 0
2
41614.3 72
0
13 SR Flip-Flop~
219 1837 372 0 4 9
0 549 497 452 496
0
0 0 4720 90
4 SRFF
-14 -53 14 -45
3 U21
25 -29 46 -21
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
12 type:digital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 0 1 0 0 0
1 U
813 0 0
2
41614.3 73
0
8 2-In OR~
219 1761 470 0 3 22
0 548 550 549
0
0 0 624 0
6 74LS32
-21 -24 21 -16
4 U12B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 8 0
1 U
3820 0 0
2
41614.3 74
0
4 4585
219 1667 485 0 14 29
0 2 554 555 556 448 449 450 451 551
552 553 548 550 608
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U19
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
3662 0 0
2
41614.3 75
0
4 4585
219 1520 346 0 14 29
0 557 558 559 560 277 459 460 461 609
495 610 553 552 551
0
0 0 4848 0
4 4585
-14 -60 14 -52
3 U18
-11 -61 10 -53
0
15 DVDD=16;DGND=8;
136 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 15 2 7 10 14 1 9 11 4
6 5 12 3 13 15 2 7 10 14
1 9 11 4 6 5 12 3 13 0
65 0 0 512 1 0 0 0
1 U
9261 0 0
2
41614.3 76
0
14 NO PushButton~
191 65 272 0 2 5
0 497 491
0
0 0 4720 0
0
5 Reset
-17 -20 18 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3447 0 0
2
41614.3 77
0
7 74LS273
150 1376 135 0 18 37
0 491 561 568 567 566 565 564 563 562
491 554 555 556 557 558 559 560 495
0
0 0 4848 0
7 74LS273
-24 -60 25 -52
3 U14
-11 -61 10 -53
0
16 DVCC=20;DGND=10;
152 %D [%20bi %10bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%20bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o %15o %16o %17o %18o] %M
0
12 type:digital
5 DIP20
37

0 1 11 18 17 14 13 8 7 4
3 19 16 15 12 9 6 5 2 1
11 18 17 14 13 8 7 4 3 19
16 15 12 9 6 5 2 0
65 0 0 0 1 0 0 0
1 U
7649 0 0
2
41614.3 78
0
8 3-In OR~
219 583 83 0 4 22
0 536 498 537 579
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 4 0
1 U
3572 0 0
2
41614.3 79
0
7 Buffer~
58 1057 611 0 2 22
0 569 546
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6F
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
9899 0 0
2
41614.3 80
0
7 Buffer~
58 850 126 0 2 22
0 587 569
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6E
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
3940 0 0
2
41614.3 81
0
12 D Flip-Flop~
219 1252 792 0 4 9
0 572 546 611 451
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U17
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
680 0 0
2
41614.3 82
0
12 D Flip-Flop~
219 1252 752 0 4 9
0 571 546 612 450
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U16
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3236 0 0
2
41614.3 83
0
12 D Flip-Flop~
219 1252 710 0 4 9
0 570 546 613 449
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U15
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5560 0 0
2
41614.3 84
0
6 74LS83
105 1008 727 0 14 29
0 448 449 450 451 511 513 573 574 575
547 570 571 572 614
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
3 U13
-10 -61 11 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 512 1 0 0 0
1 U
3609 0 0
2
41614.3 85
0
7 Buffer~
58 553 683 0 2 22
0 576 574
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6D
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
4752 0 0
2
41614.3 86
0
7 Buffer~
58 552 643 0 2 22
0 577 573
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6C
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
6635 0 0
2
41614.3 87
0
9 2-In AND~
219 495 585 0 3 22
0 581 580 577
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11B
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 7 0
1 U
5511 0 0
2
41614.3 88
0
9 Inverter~
13 510 531 0 2 22
0 580 581
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3F
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
7227 0 0
2
41614.3 89
0
9 2-In AND~
219 432 583 0 3 22
0 582 545 576
0
0 0 624 270
6 74LS08
-21 -24 21 -16
4 U11A
13 -4 41 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
8673 0 0
2
41614.3 90
0
9 Inverter~
13 447 529 0 2 22
0 545 582
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3E
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
5175 0 0
2
41614.3 91
0
8 2-In OR~
219 682 66 0 3 22
0 578 579 561
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U5B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 6 0
1 U
9215 0 0
2
41614.3 92
0
8 3-In OR~
219 585 44 0 4 22
0 539 538 541 578
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
3186 0 0
2
41614.3 93
0
14 NO PushButton~
191 63 226 0 2 5
0 537 491
0
0 0 4720 0
0
7 HalfDol
-25 -20 24 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3894 0 0
2
41614.3 94
0
14 NO PushButton~
191 62 179 0 2 5
0 536 491
0
0 0 4720 0
0
7 Quarter
-24 -20 25 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3898 0 0
2
41614.3 95
0
14 NO PushButton~
191 66 131 0 2 5
0 541 491
0
0 0 4720 0
0
4 Dime
-14 -20 14 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
362 0 0
2
41614.3 96
0
14 NO PushButton~
191 68 91 0 2 5
0 538 491
0
0 0 4720 0
0
6 Nickle
-21 -20 21 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
3755 0 0
2
41614.3 97
0
14 NO PushButton~
191 73 44 0 2 5
0 539 491
0
0 0 4720 0
0
5 Penny
-17 -20 18 -12
0
0
0
0
0
4 SIP2
5

0 1 2 1 2 0
0 0 0 0 1 0 0 0
1 S
4103 0 0
2
41614.3 98
0
7 Ground~
168 34 787 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3992 0 0
2
41614.3 99
0
2 +V
167 13 16 0 1 3
0 491
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4205 0 0
2
41614.3 100
0
12 D Flip-Flop~
219 1057 440 0 4 9
0 586 569 615 461
0
0 0 4720 0
3 DFF
-10 -53 11 -45
3 U10
-11 -55 10 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
5841 0 0
2
5.89641e-315 5.56337e-315
0
12 D Flip-Flop~
219 1055 396 0 4 9
0 585 569 616 460
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U9
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
8703 0 0
2
5.89641e-315 5.5637e-315
0
12 D Flip-Flop~
219 1053 353 0 4 9
0 584 569 617 459
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U8
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
4198 0 0
2
5.89641e-315 5.56402e-315
0
12 D Flip-Flop~
219 1052 307 0 4 9
0 583 569 618 277
0
0 0 4720 0
3 DFF
-10 -53 11 -45
2 U7
-7 -55 7 -47
0
14 DVCC=6;DGND=5;
47 %D [%6bi %5bi %1i %2i][%6bo %1o %2o %3o %4o] %M
0
11 typeDigital
4 DIP6
9

0 1 2 3 4 1 2 3 4 0
65 0 0 512 1 0 0 0
1 U
3495 0 0
2
5.89641e-315 5.56435e-315
0
7 Buffer~
58 818 169 0 2 22
0 561 587
0
0 0 624 0
4 4050
-14 -19 14 -11
3 U6B
-11 -20 10 -12
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
5247 0 0
2
5.89641e-315 5.56467e-315
0
9 Inverter~
13 404 278 0 2 22
0 542 592
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3D
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
3399 0 0
2
5.89641e-315 5.56499e-315
0
9 2-In AND~
219 389 332 0 3 22
0 592 542 591
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 3 0
1 U
7916 0 0
2
5.89641e-315 5.56532e-315
0
9 Inverter~
13 330 278 0 2 22
0 544 593
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3C
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3913 0 0
2
5.89641e-315 5.56564e-315
0
9 2-In AND~
219 315 332 0 3 22
0 593 544 590
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 3 0
1 U
729 0 0
2
5.89641e-315 5.56596e-315
0
9 Inverter~
13 258 280 0 2 22
0 543 594
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
3882 0 0
2
5.89641e-315 5.56629e-315
0
9 2-In AND~
219 243 334 0 3 22
0 594 543 589
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
5428 0 0
2
5.89641e-315 5.56661e-315
0
9 2-In AND~
219 181 325 0 3 22
0 595 540 588
0
0 0 624 270
6 74LS08
-21 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
6908 0 0
2
5.89641e-315 5.56694e-315
0
9 Inverter~
13 196 271 0 2 22
0 540 595
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U3A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
5761 0 0
2
5.89641e-315 5.56726e-315
0
6 74LS83
105 869 375 0 14 29
0 277 459 460 461 591 590 589 588 2
583 584 585 586 575
0
0 0 4848 0
6 74LS83
-21 -60 21 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3416 0 0
2
5.89641e-315 5.56758e-315
0
9 Resistor~
219 249 511 0 3 5
0 2 497 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R6
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 22
82 0 0 0 1 0 0 0
1 R
3390 0 0
2
41614.3 101
0
9 Resistor~
219 210 511 0 3 5
0 2 537 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 26
82 0 0 0 1 0 0 0
1 R
3425 0 0
2
41614.3 102
0
9 Resistor~
219 178 513 0 3 5
0 2 536 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
692 0 0
2
41614.3 103
0
9 Resistor~
219 147 512 0 3 5
0 2 541 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 62
82 0 0 0 1 0 0 0
1 R
5714 0 0
2
41614.3 104
0
9 Resistor~
219 116 512 0 3 5
0 2 538 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 106
82 0 0 0 1 0 0 0
1 R
354 0 0
2
41614.3 105
0
9 Resistor~
219 80 511 0 3 5
0 2 539 -1
0
0 0 880 90
2 1k
8 0 22 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 50
82 0 0 0 1 0 0 0
1 R
9446 0 0
2
41614.3 106
0
982
0 0 3 0 0 4096 0 0 0 11 36 3
1247 3450
1304 3450
1304 3416
1 0 3 0 0 12288 0 16 0 0 11 4
618 2168
634 2168
634 2134
709 2134
0 1 3 0 0 16 0 0 9 11 0 2
709 2062
649 2062
2 0 4 0 0 4112 0 8 0 0 352 3
576 2030
658 2030
658 2009
3 0 5 0 0 8208 0 8 0 0 26 3
531 2039
504 2039
504 2009
1 2 6 0 0 4240 0 8 9 0 0 4
576 2048
605 2048
605 2062
613 2062
0 1 3 0 0 4096 0 0 15 11 0 2
709 1945
613 1945
1 0 3 0 0 0 0 14 0 0 11 4
613 1876
704 1876
704 1877
709 1877
0 1 3 0 0 0 0 0 10 11 0 2
709 1774
648 1774
0 1 3 0 0 4096 0 0 13 11 0 2
709 1678
610 1678
0 1 3 0 0 12416 0 0 12 0 0 5
1247 3419
1247 3471
709 3471
709 1603
610 1603
2 0 7 0 0 4096 0 16 0 0 351 3
618 2150
663 2150
663 2122
3 0 8 0 0 8192 0 16 0 0 25 3
572 2159
549 2159
549 2122
3 0 9 0 0 4096 0 15 0 0 27 3
567 1936
537 1936
537 1907
2 0 10 0 0 4096 0 15 0 0 353 3
613 1927
661 1927
661 1907
2 0 11 0 0 4096 0 14 0 0 354 3
613 1858
660 1858
660 1841
2 0 12 0 0 4096 0 11 0 0 373 3
575 1742
657 1742
657 1718
3 0 13 0 0 8192 0 11 0 0 29 3
530 1751
503 1751
503 1718
3 0 14 0 0 4096 0 14 0 0 28 3
567 1867
539 1867
539 1841
2 0 15 0 0 4096 0 13 0 0 374 3
610 1660
663 1660
663 1646
3 0 16 0 0 4096 0 13 0 0 30 3
564 1669
537 1669
537 1646
2 0 17 0 0 4096 0 12 0 0 375 3
610 1585
659 1585
659 1571
0 3 18 0 0 8192 0 0 12 31 0 3
526 1571
526 1594
564 1594
1 2 19 0 0 4224 0 11 10 0 0 4
575 1760
604 1760
604 1774
612 1774
0 0 8 0 0 4096 0 0 0 0 725 2
597 2122
453 2122
0 0 5 0 0 4096 0 0 0 0 726 2
600 2009
440 2009
0 0 9 0 0 4096 0 0 0 0 727 2
601 1907
433 1907
0 0 14 0 0 4096 0 0 0 0 728 2
606 1841
423 1841
0 0 13 0 0 4096 0 0 0 0 729 2
600 1718
411 1718
0 0 16 0 0 4096 0 0 0 0 730 2
601 1646
406 1646
0 0 18 0 0 4096 0 0 0 0 731 2
590 1571
399 1571
1 0 3 0 0 0 0 19 0 0 36 2
1143 3229
1567 3229
1 0 3 0 0 0 0 20 0 0 36 2
1145 3269
1567 3269
1 0 3 0 0 0 0 21 0 0 36 2
1152 3313
1567 3313
1 0 3 0 0 0 0 22 0 0 36 2
1159 3360
1567 3360
0 1 3 0 0 0 0 0 23 37 0 3
1567 3155
1567 3416
1163 3416
0 1 3 0 0 0 0 0 17 594 0 5
2356 2739
2356 3053
1643 3053
1643 3155
1136 3155
2 0 20 0 0 4096 0 17 0 0 113 3
1136 3137
1194 3137
1194 3131
2 0 21 0 0 4096 0 18 0 0 112 3
1140 3177
1193 3177
1193 3169
2 0 22 0 0 4096 0 19 0 0 111 3
1143 3211
1199 3211
1199 3204
2 0 23 0 0 4096 0 20 0 0 110 3
1145 3251
1201 3251
1201 3241
2 0 24 0 0 4096 0 21 0 0 109 3
1152 3295
1204 3295
1204 3282
2 0 25 0 0 4096 0 22 0 0 108 3
1159 3342
1209 3342
1209 3328
2 0 26 0 0 4096 0 23 0 0 107 3
1163 3398
1206 3398
1206 3375
3 0 27 0 0 8192 0 23 0 0 52 3
1117 3407
1086 3407
1086 3375
3 0 28 0 0 4096 0 22 0 0 53 3
1113 3351
1089 3351
1089 3328
3 0 29 0 0 8192 0 21 0 0 54 3
1106 3304
1086 3304
1086 3282
3 0 30 0 0 8192 0 20 0 0 55 3
1099 3260
1081 3260
1081 3241
3 0 31 0 0 4096 0 19 0 0 56 3
1097 3220
1079 3220
1079 3204
3 0 32 0 0 8192 0 18 0 0 57 3
1094 3186
1083 3186
1083 3169
3 0 33 0 0 8192 0 17 0 0 58 3
1090 3146
1076 3146
1076 3131
0 0 27 0 0 8192 0 0 0 0 657 4
1144 3375
924 3375
924 2221
775 2221
0 0 28 0 0 8192 0 0 0 0 658 6
1137 3328
947 3328
947 2286
903 2286
903 2210
765 2210
0 0 29 0 0 16384 0 0 0 0 659 6
1124 3282
1001 3282
1001 2813
960 2813
960 2200
755 2200
0 0 30 0 0 8192 0 0 0 0 660 4
1123 3241
697 3241
697 2190
745 2190
0 0 31 0 0 8192 0 0 0 0 661 4
1117 3204
679 3204
679 2176
735 2176
0 0 32 0 0 8192 0 0 0 0 662 4
1109 3169
661 3169
661 2167
725 2167
0 0 33 0 0 8192 0 0 0 0 663 4
1094 3131
647 3131
647 2157
792 2157
2 1 34 0 0 12416 0 24 80 0 0 4
3263 3029
3263 3038
3256 3038
3256 3053
4 1 35 0 0 4224 0 25 24 0 0 4
3269 2977
3269 2985
3263 2985
3263 2993
2 1 36 0 0 4224 0 27 82 0 0 4
3173 3032
3173 3041
3166 3041
3166 3049
2 2 37 0 0 12416 0 26 80 0 0 4
3233 3030
3233 3038
3238 3038
3238 3053
4 1 38 0 0 4224 0 31 26 0 0 4
3229 2974
3229 2986
3233 2986
3233 2994
4 1 39 0 0 4224 0 32 27 0 0 4
3174 2975
3174 2988
3173 2988
3173 2996
2 1 40 0 0 4224 0 28 84 0 0 3
3089 3030
3089 3043
3077 3043
4 1 41 0 0 12416 0 33 28 0 0 4
3087 2979
3087 2986
3089 2986
3089 2994
2 1 42 0 0 8320 0 29 86 0 0 3
2998 3028
2998 3040
2985 3040
4 1 43 0 0 12416 0 34 29 0 0 4
2999 2979
2999 2984
2998 2984
2998 2992
2 1 44 0 0 8320 0 30 87 0 0 3
2909 3028
2909 3038
2898 3038
4 1 45 0 0 4224 0 35 30 0 0 2
2909 2976
2909 2992
3 0 46 0 0 4096 0 35 0 0 239 2
2900 2931
2899 2931
2 0 47 0 0 4096 0 35 0 0 238 2
2909 2931
2908 2931
1 0 48 0 0 4096 0 35 0 0 237 2
2918 2931
2917 2931
2 1 49 0 0 4224 0 37 90 0 0 3
2729 3022
2729 3037
2721 3037
2 1 50 0 0 8320 0 38 91 0 0 4
2653 3018
2653 3022
2637 3022
2637 3034
2 1 51 0 0 4224 0 39 122 0 0 3
2560 3017
2560 3029
2549 3029
2 1 52 0 0 8320 0 36 89 0 0 3
2823 3023
2823 3037
2806 3037
4 1 53 0 0 8320 0 40 36 0 0 4
2815 2975
2815 2979
2823 2979
2823 2987
4 1 54 0 0 4224 0 41 37 0 0 3
2730 2977
2730 2986
2729 2986
4 1 55 0 0 4224 0 42 38 0 0 3
2650 2975
2650 2982
2653 2982
4 1 56 0 0 12416 0 43 39 0 0 4
2559 2970
2559 2975
2560 2975
2560 2981
2 2 57 0 0 4224 0 44 89 0 0 3
2779 3023
2779 3037
2788 3037
4 1 58 0 0 12416 0 48 44 0 0 4
2776 2975
2776 2979
2779 2979
2779 2987
2 2 59 0 0 4224 0 45 90 0 0 3
2690 3024
2690 3037
2703 3037
4 1 60 0 0 12416 0 49 45 0 0 4
2692 2974
2692 2980
2690 2980
2690 2988
2 2 61 0 0 8320 0 46 91 0 0 4
2607 3018
2607 3022
2619 3022
2619 3034
4 1 62 0 0 4224 0 50 46 0 0 2
2607 2971
2607 2982
2 2 63 0 0 4224 0 47 122 0 0 3
2523 3015
2523 3029
2531 3029
4 1 64 0 0 12416 0 51 47 0 0 4
2520 2968
2520 2973
2523 2973
2523 2979
3 0 65 0 0 0 0 50 0 0 262 2
2598 2926
2598 2926
2 0 66 0 0 0 0 50 0 0 261 2
2607 2926
2607 2926
1 0 67 0 0 0 0 50 0 0 260 2
2616 2926
2616 2926
1 4 68 0 0 4224 0 54 57 0 0 4
2502 283
2502 301
2508 301
2508 308
1 4 69 0 0 4224 0 53 56 0 0 4
2732 275
2732 293
2738 293
2738 300
1 4 70 0 0 4224 0 52 55 0 0 4
2839 277
2839 291
2846 291
2846 298
2 2 71 0 0 4224 0 52 111 0 0 4
2839 241
2839 225
2827 225
2827 210
2 2 72 0 0 12416 0 53 113 0 0 4
2732 239
2732 227
2726 227
2726 212
2 2 73 0 0 4224 0 54 116 0 0 4
2502 247
2502 229
2494 229
2494 214
3 0 74 0 0 4096 0 57 0 0 336 2
2517 353
2518 353
2 0 75 0 0 4096 0 57 0 0 337 2
2508 353
2509 353
1 0 76 0 0 4096 0 57 0 0 338 2
2499 353
2500 353
1 4 77 0 0 4224 0 58 59 0 0 4
2630 272
2630 293
2636 293
2636 300
2 2 78 0 0 4224 0 115 58 0 0 4
2620 212
2620 228
2630 228
2630 236
4 0 79 0 0 4096 0 119 0 0 191 2
3066 1103
3066 1212
0 3 80 0 0 4096 0 0 93 141 0 2
3368 187
3368 226
2 0 81 0 0 4096 0 62 0 0 128 2
1725 3286
1820 3286
4 0 26 0 0 4224 0 61 0 0 0 2
1674 3375
1148 3375
5 0 25 0 0 4224 0 63 0 0 0 2
1670 3328
1141 3328
5 0 24 0 0 4224 0 62 0 0 0 2
1675 3282
1128 3282
4 0 23 0 0 4224 0 60 0 0 0 2
1671 3241
1127 3241
2 0 22 0 0 4224 0 64 0 0 0 2
1681 3204
1121 3204
3 0 21 0 0 4224 0 65 0 0 0 2
1669 3169
1113 3169
3 0 20 0 0 4224 0 66 0 0 0 2
1667 3131
1098 3131
1 0 82 0 0 4096 0 61 0 0 124 3
1726 3384
1869 3384
1869 3370
2 0 83 0 0 8320 0 61 0 0 131 3
1725 3375
1839 3375
1839 3122
3 0 84 0 0 8320 0 61 0 0 123 3
1726 3366
1827 3366
1827 3088
0 2 82 0 0 8192 0 0 63 124 0 4
1897 3370
1897 3336
1726 3336
1726 3332
3 1 85 0 0 8320 0 73 63 0 0 4
1920 3210
1856 3210
1856 3341
1726 3341
3 0 86 0 0 8192 0 63 0 0 127 3
1726 3323
1876 3323
1876 3167
4 0 83 0 0 0 0 63 0 0 131 3
1726 3314
1886 3314
1886 3122
3 1 87 0 0 8320 0 68 62 0 0 4
1919 3411
1809 3411
1809 3295
1725 3295
0 3 86 0 0 8320 0 0 62 127 0 3
1891 3167
1891 3277
1725 3277
3 4 84 0 0 0 0 76 62 0 0 4
1921 3088
1789 3088
1789 3268
1725 3268
3 1 82 0 0 4224 0 69 60 0 0 4
1917 3370
1745 3370
1745 3250
1723 3250
2 0 88 0 0 4096 0 60 0 0 130 2
1722 3241
1836 3241
0 3 83 0 0 0 0 0 60 131 0 3
1866 3122
1866 3232
1723 3232
1 3 86 0 0 0 0 64 74 0 0 4
1717 3204
1863 3204
1863 3167
1920 3167
1 3 81 0 0 8320 0 65 70 0 0 4
1721 3178
1820 3178
1820 3331
1919 3331
2 3 89 0 0 8320 0 65 71 0 0 4
1721 3160
1829 3160
1829 3290
1919 3290
1 3 88 0 0 4224 0 66 72 0 0 4
1719 3140
1836 3140
1836 3249
1919 3249
2 3 83 0 0 0 0 66 75 0 0 4
1719 3122
1929 3122
1929 3126
1923 3126
3 1 90 0 0 12416 0 116 76 0 0 5
2485 168
2485 94
3457 94
3457 3097
1967 3097
3 1 91 0 0 12416 0 115 75 0 0 5
2611 166
2611 100
3463 100
3463 3135
1969 3135
3 1 92 0 0 12416 0 113 74 0 0 5
2717 166
2717 107
3470 107
3470 3176
1966 3176
3 1 93 0 0 12416 0 111 73 0 0 5
2818 164
2818 116
3477 116
3477 3219
1966 3219
3 1 94 0 0 12416 0 108 72 0 0 5
2912 227
2912 124
3484 124
3484 3258
1965 3258
3 1 95 0 0 12416 0 105 71 0 0 5
3002 225
3002 136
3493 136
3493 3299
1965 3299
3 1 96 0 0 12416 0 102 70 0 0 5
3091 223
3091 150
3503 150
3503 3340
1965 3340
3 1 97 0 0 12416 0 99 69 0 0 5
3184 223
3184 163
3519 163
3519 3379
1963 3379
3 1 98 0 0 12416 0 96 68 0 0 5
3277 224
3277 176
3533 176
3533 3420
1965 3420
0 1 80 0 0 12416 0 0 67 0 0 5
3367 233
3367 187
3546 187
3546 3456
1965 3456
3 2 99 0 0 8320 0 79 67 0 0 3
3336 3041
3336 3438
1965 3438
3 2 100 0 0 8320 0 80 68 0 0 3
3247 3099
3247 3402
1965 3402
3 2 101 0 0 8320 0 82 69 0 0 3
3157 3095
3157 3361
1963 3361
3 2 102 0 0 8320 0 84 70 0 0 3
3068 3089
3068 3322
1965 3322
3 2 103 0 0 8320 0 86 71 0 0 3
2976 3086
2976 3281
1965 3281
3 2 104 0 0 8320 0 87 72 0 0 3
2889 3084
2889 3240
1965 3240
3 2 105 0 0 8320 0 89 73 0 0 3
2797 3083
2797 3201
1966 3201
3 2 106 0 0 8320 0 90 74 0 0 3
2712 3083
2712 3158
1966 3158
3 2 107 0 0 8320 0 91 75 0 0 3
2628 3080
2628 3117
1969 3117
3 2 108 0 0 8320 0 122 76 0 0 3
2540 3075
2540 3079
1967 3079
2 0 109 0 0 4096 0 124 0 0 153 2
3398 2161
3398 2133
0 1 109 0 0 8320 0 0 124 350 0 4
1723 2753
1723 2133
3407 2133
3407 2161
2 0 110 0 0 4096 0 123 0 0 155 2
3251 2160
3251 2137
0 1 110 0 0 8320 0 0 123 603 0 4
1723 2536
1723 2137
3260 2137
3260 2160
2 0 111 0 0 4096 0 125 0 0 157 2
3105 2160
3105 2142
0 1 111 0 0 8320 0 0 125 605 0 4
1726 2371
1726 2142
3114 2142
3114 2160
0 2 112 0 0 4096 0 0 126 159 0 2
2955 2147
2955 2160
0 1 112 0 0 8320 0 0 126 607 0 4
1721 2208
1721 2147
2964 2147
2964 2160
2 0 113 0 0 4096 0 121 0 0 161 2
3395 1110
3395 1133
0 1 113 0 0 8320 0 0 121 609 0 4
1716 2040
1716 1133
3404 1133
3404 1110
1 0 114 0 0 8192 0 120 0 0 163 4
3257 1109
3257 1122
3239 1122
3239 1127
0 2 114 0 0 8320 0 0 120 611 0 4
1714 1877
1714 1127
3248 1127
3248 1109
0 2 115 0 0 4096 0 0 119 165 0 2
3102 1122
3102 1109
0 1 115 0 0 8320 0 0 119 613 0 4
1714 1772
1714 1122
3111 1122
3111 1109
0 1 116 0 0 4096 0 0 118 167 0 3
2952 1117
2961 1117
2961 1109
0 2 116 0 0 8320 0 0 118 615 0 4
1701 1608
1701 1117
2952 1117
2952 1109
6 0 117 0 0 4096 0 125 0 0 170 2
3051 2166
3051 2121
6 0 117 0 0 0 0 123 0 0 170 2
3197 2166
3197 2121
0 6 117 0 0 4096 0 0 124 180 0 3
2894 2121
3344 2121
3344 2167
5 0 118 0 0 4096 0 125 0 0 173 2
3060 2166
3060 2111
5 0 118 0 0 0 0 123 0 0 173 2
3206 2166
3206 2111
0 5 118 0 0 4096 0 0 124 181 0 3
2910 2111
3353 2111
3353 2167
4 0 79 0 0 0 0 125 0 0 176 2
3069 2166
3069 2103
4 0 79 0 0 0 0 123 0 0 176 2
3215 2166
3215 2103
0 4 79 0 0 4096 0 0 124 182 0 3
2914 2103
3362 2103
3362 2167
3 0 119 0 0 4096 0 125 0 0 179 2
3078 2166
3078 2097
3 0 119 0 0 0 0 123 0 0 179 2
3224 2166
3224 2097
0 3 119 0 0 4096 0 0 124 183 0 3
2923 2097
3371 2097
3371 2167
0 6 117 0 0 4096 0 0 126 198 0 4
2894 1187
2894 2152
2901 2152
2901 2166
0 5 118 0 0 8192 0 0 126 197 0 3
2907 1211
2910 1211
2910 2166
0 4 79 0 0 4096 0 0 126 196 0 4
2914 1237
2914 2152
2919 2152
2919 2166
0 3 119 0 0 4096 0 0 126 195 0 4
2923 1262
2923 2152
2928 2152
2928 2166
6 0 117 0 0 0 0 119 0 0 186 2
3048 1103
3048 1175
6 0 117 0 0 0 0 120 0 0 186 2
3194 1103
3194 1175
0 6 117 0 0 0 0 0 121 198 0 3
2898 1175
3341 1175
3341 1104
5 0 118 0 0 0 0 119 0 0 189 2
3057 1103
3057 1194
5 0 118 0 0 0 0 120 0 0 189 2
3203 1103
3203 1194
0 5 118 0 0 0 0 0 121 197 0 3
2907 1194
3350 1194
3350 1104
4 0 79 0 0 0 0 120 0 0 191 2
3212 1103
3212 1212
0 4 79 0 0 0 0 0 121 196 0 3
2916 1212
3359 1212
3359 1104
3 0 119 0 0 0 0 119 0 0 194 2
3075 1103
3075 1232
3 0 119 0 0 0 0 120 0 0 194 2
3221 1103
3221 1232
0 3 119 0 0 0 0 0 121 195 0 5
2925 1232
3369 1232
3369 1092
3368 1092
3368 1104
0 3 119 0 0 0 0 0 118 672 0 3
2412 1262
2925 1262
2925 1103
0 4 79 0 0 0 0 0 118 674 0 3
2302 1237
2916 1237
2916 1103
0 5 118 0 0 0 0 0 118 676 0 3
2194 1215
2907 1215
2907 1103
0 6 117 0 0 0 0 0 118 678 0 3
2074 1187
2898 1187
2898 1103
1 15 120 0 0 4224 0 78 124 0 0 4
3364 2931
3364 2250
3380 2250
3380 2237
2 9 121 0 0 4224 0 78 123 0 0 4
3355 2931
3355 2269
3287 2269
3287 2236
3 19 122 0 0 4224 0 78 123 0 0 4
3346 2931
3346 2314
3197 2314
3197 2236
1 13 123 0 0 4224 0 77 125 0 0 4
3325 2929
3325 2374
3105 2374
3105 2236
2 7 124 0 0 4224 0 77 126 0 0 4
3316 2929
3316 2404
3009 2404
3009 2236
3 17 125 0 0 4224 0 77 126 0 0 4
3307 2929
3307 2399
2919 2399
2919 2236
1 16 126 0 0 8320 0 25 124 0 0 5
3278 2932
3277 2932
3277 2245
3371 2245
3371 2237
2 10 127 0 0 8320 0 25 123 0 0 5
3269 2932
3268 2932
3268 2269
3278 2269
3278 2236
3 20 128 0 0 8320 0 25 123 0 0 5
3260 2932
3259 2932
3259 2289
3188 2289
3188 2236
1 14 129 0 0 4224 0 31 125 0 0 4
3238 2929
3238 2369
3096 2369
3096 2236
2 8 130 0 0 4224 0 31 126 0 0 4
3229 2929
3229 2394
3000 2394
3000 2236
3 18 131 0 0 4224 0 31 126 0 0 4
3220 2929
3220 2389
2910 2389
2910 2236
4 1 132 0 0 4224 0 78 79 0 0 3
3355 2982
3355 2995
3345 2995
4 2 133 0 0 4224 0 77 79 0 0 3
3316 2980
3316 2995
3327 2995
1 7 134 0 0 4224 0 32 124 0 0 4
3183 2930
3183 2265
3452 2265
3452 2237
2 17 135 0 0 4224 0 32 124 0 0 4
3174 2930
3174 2285
3362 2285
3362 2237
3 11 136 0 0 4224 0 32 123 0 0 4
3165 2930
3165 2244
3269 2244
3269 2236
1 21 137 0 0 4224 0 81 123 0 0 4
3150 2932
3150 2264
3179 2264
3179 2236
3 15 138 0 0 4224 0 81 125 0 0 4
3138 2932
3138 2344
3087 2344
3087 2236
2 9 139 0 0 4224 0 81 126 0 0 4
3126 2932
3126 2384
2991 2384
2991 2236
4 19 140 0 0 4224 0 81 126 0 0 4
3114 2932
3114 2379
2901 2379
2901 2236
1 8 141 0 0 4224 0 33 124 0 0 4
3096 2934
3096 2310
3443 2310
3443 2237
2 18 142 0 0 4224 0 33 124 0 0 4
3087 2934
3087 2250
3353 2250
3353 2237
3 12 143 0 0 4224 0 33 123 0 0 4
3078 2934
3078 2279
3260 2279
3260 2236
1 22 144 0 0 4224 0 83 123 0 0 4
3063 2935
3063 2284
3170 2284
3170 2236
3 16 145 0 0 4224 0 83 125 0 0 4
3051 2935
3051 2249
3078 2249
3078 2236
2 10 146 0 0 4224 0 83 126 0 0 4
3039 2935
3039 2374
2982 2374
2982 2236
4 20 147 0 0 4224 0 83 126 0 0 4
3027 2935
3027 2369
2892 2369
2892 2236
1 9 148 0 0 8320 0 34 124 0 0 5
3008 2934
3007 2934
3007 2365
3434 2365
3434 2237
2 19 149 0 0 8320 0 34 124 0 0 5
2999 2934
2998 2934
2998 2340
3344 2340
3344 2237
3 13 150 0 0 8320 0 34 123 0 0 5
2990 2934
2989 2934
2989 2304
3251 2304
3251 2236
1 7 151 0 0 4224 0 85 125 0 0 4
2974 2936
2974 2244
3159 2244
3159 2236
3 17 152 0 0 4224 0 85 125 0 0 4
2962 2936
2962 2279
3069 2279
3069 2236
2 11 153 0 0 4224 0 85 126 0 0 4
2950 2936
2950 2244
2973 2244
2973 2236
4 21 154 0 0 4224 0 85 126 0 0 4
2938 2936
2938 2364
2883 2364
2883 2236
5 2 155 0 0 12416 0 81 82 0 0 4
3132 2983
3132 2989
3148 2989
3148 3049
5 2 156 0 0 12416 0 83 84 0 0 4
3045 2986
3045 2992
3059 2992
3059 3043
5 2 157 0 0 12416 0 85 86 0 0 4
2956 2987
2956 2993
2967 2993
2967 3040
0 10 48 0 0 4224 0 0 124 0 0 4
2917 2935
2917 2360
3425 2360
3425 2237
0 20 47 0 0 4224 0 0 124 0 0 4
2908 2935
2908 2355
3335 2355
3335 2237
0 14 46 0 0 4224 0 0 123 0 0 4
2899 2935
2899 2349
3242 2349
3242 2236
1 8 158 0 0 4224 0 88 125 0 0 4
2884 2935
2884 2334
3150 2334
3150 2236
3 18 159 0 0 4224 0 88 125 0 0 4
2872 2935
2872 2344
3060 2344
3060 2236
2 12 160 0 0 4224 0 88 126 0 0 4
2860 2935
2860 2339
2964 2339
2964 2236
4 22 161 0 0 4224 0 88 126 0 0 4
2848 2935
2848 2334
2874 2334
2874 2236
5 2 162 0 0 12416 0 88 87 0 0 4
2866 2986
2866 2992
2880 2992
2880 3038
1 11 163 0 0 4224 0 40 124 0 0 4
2824 2930
2824 2330
3416 2330
3416 2237
2 21 164 0 0 4224 0 40 124 0 0 4
2815 2930
2815 2325
3326 2325
3326 2237
3 15 165 0 0 4224 0 40 123 0 0 4
2806 2930
2806 2319
3233 2319
3233 2236
1 9 166 0 0 4224 0 48 125 0 0 4
2785 2930
2785 2314
3141 2314
3141 2236
2 19 167 0 0 4224 0 48 125 0 0 4
2776 2930
2776 2309
3051 2309
3051 2236
3 13 168 0 0 4224 0 48 126 0 0 4
2767 2930
2767 2304
2955 2304
2955 2236
1 12 169 0 0 4224 0 41 124 0 0 4
2739 2932
2739 2260
3407 2260
3407 2237
2 22 170 0 0 4224 0 41 124 0 0 4
2730 2932
2730 2300
3317 2300
3317 2237
3 16 171 0 0 4224 0 41 123 0 0 4
2721 2932
2721 2294
3224 2294
3224 2236
1 10 172 0 0 8320 0 49 125 0 0 5
2701 2929
2700 2929
2700 2289
3132 2289
3132 2236
2 20 173 0 0 8320 0 49 125 0 0 5
2692 2929
2691 2929
2691 2284
3042 2284
3042 2236
3 14 174 0 0 8320 0 49 126 0 0 5
2683 2929
2682 2929
2682 2279
2946 2279
2946 2236
1 13 175 0 0 8320 0 42 124 0 0 4
2659 2930
2659 2255
3398 2255
3398 2237
2 7 176 0 0 4224 0 42 123 0 0 4
2650 2930
2650 2274
3305 2274
3305 2236
3 17 177 0 0 4224 0 42 123 0 0 4
2641 2930
2641 2269
3215 2269
3215 2236
0 11 67 0 0 4224 0 0 125 0 0 4
2616 2930
2616 2264
3123 2264
3123 2236
0 21 66 0 0 4224 0 0 125 0 0 4
2607 2930
2607 2249
3033 2249
3033 2236
0 15 65 0 0 4224 0 0 126 0 0 4
2598 2930
2598 2244
2937 2244
2937 2236
2 11 178 0 0 4224 0 94 121 0 0 4
3400 342
3400 1021
3413 1021
3413 1034
1 21 179 0 0 4224 0 94 121 0 0 4
3382 342
3382 1021
3323 1021
3323 1034
4 15 180 0 0 4224 0 92 120 0 0 4
3361 342
3361 980
3230 980
3230 1033
2 9 181 0 0 4224 0 92 119 0 0 4
3349 342
3349 940
3138 940
3138 1033
3 19 182 0 0 4224 0 92 119 0 0 4
3337 342
3337 945
3048 945
3048 1033
1 13 183 0 0 4224 0 92 118 0 0 4
3325 342
3325 950
2952 950
2952 1033
2 12 184 0 0 4224 0 97 121 0 0 4
3309 340
3309 1026
3404 1026
3404 1034
1 22 185 0 0 4224 0 97 121 0 0 4
3291 340
3291 1011
3314 1011
3314 1034
4 16 186 0 0 4224 0 95 120 0 0 4
3270 340
3270 985
3221 985
3221 1033
2 10 187 0 0 4224 0 95 119 0 0 4
3258 340
3258 955
3129 955
3129 1033
3 20 188 0 0 4224 0 95 119 0 0 4
3246 340
3246 960
3039 960
3039 1033
1 14 189 0 0 4224 0 95 118 0 0 4
3234 340
3234 965
2943 965
2943 1033
2 13 190 0 0 4224 0 100 121 0 0 4
3216 339
3216 1016
3395 1016
3395 1034
1 7 191 0 0 4224 0 100 120 0 0 4
3198 339
3198 1025
3302 1025
3302 1033
4 17 192 0 0 4224 0 98 120 0 0 4
3177 339
3177 980
3212 980
3212 1033
2 11 193 0 0 4224 0 98 119 0 0 4
3165 339
3165 970
3120 970
3120 1033
3 21 194 0 0 4224 0 98 119 0 0 4
3153 339
3153 975
3030 975
3030 1033
1 15 195 0 0 4224 0 98 118 0 0 4
3141 339
3141 980
2934 980
2934 1033
2 14 196 0 0 4224 0 103 121 0 0 4
3123 339
3123 991
3386 991
3386 1034
1 8 197 0 0 4224 0 103 120 0 0 4
3105 339
3105 1020
3293 1020
3293 1033
4 18 198 0 0 4224 0 101 120 0 0 4
3084 339
3084 985
3203 985
3203 1033
2 12 199 0 0 4224 0 101 119 0 0 4
3072 339
3072 990
3111 990
3111 1033
3 22 200 0 0 4224 0 101 119 0 0 4
3060 339
3060 985
3021 985
3021 1033
1 16 201 0 0 4224 0 101 118 0 0 4
3048 339
3048 990
2925 990
2925 1033
2 15 202 0 0 4224 0 106 121 0 0 4
3034 341
3034 996
3377 996
3377 1034
1 9 203 0 0 4224 0 106 120 0 0 4
3016 341
3016 1000
3284 1000
3284 1033
4 19 204 0 0 4224 0 104 120 0 0 4
2995 341
2995 1015
3194 1015
3194 1033
2 13 205 0 0 4224 0 104 119 0 0 4
2983 341
2983 1020
3102 1020
3102 1033
3 7 206 0 0 4224 0 104 118 0 0 4
2971 341
2971 1000
3006 1000
3006 1033
1 17 207 0 0 4224 0 104 118 0 0 4
2959 341
2959 1000
2916 1000
2916 1033
3 2 208 0 0 12416 0 94 93 0 0 5
3391 291
3392 291
3392 287
3377 287
3377 272
5 1 209 0 0 8320 0 92 93 0 0 4
3343 291
3343 287
3359 287
3359 272
3 2 210 0 0 12416 0 97 96 0 0 5
3300 289
3301 289
3301 285
3286 285
3286 270
5 1 211 0 0 8320 0 95 96 0 0 4
3252 289
3252 285
3268 285
3268 270
3 2 212 0 0 12416 0 100 99 0 0 5
3207 288
3208 288
3208 284
3193 284
3193 269
5 1 213 0 0 8320 0 98 99 0 0 4
3159 288
3159 284
3175 284
3175 269
3 2 214 0 0 12416 0 103 102 0 0 5
3114 288
3115 288
3115 284
3100 284
3100 269
5 1 215 0 0 8320 0 101 102 0 0 4
3066 288
3066 284
3082 284
3082 269
3 2 216 0 0 12416 0 106 105 0 0 5
3025 290
3026 290
3026 286
3011 286
3011 271
5 1 217 0 0 8320 0 104 105 0 0 4
2977 290
2977 286
2993 286
2993 271
2 16 218 0 0 4224 0 107 121 0 0 4
2944 343
2944 1006
3368 1006
3368 1034
1 10 219 0 0 4224 0 107 120 0 0 4
2926 343
2926 1010
3275 1010
3275 1033
4 20 220 0 0 4224 0 109 120 0 0 4
2905 343
2905 1025
3185 1025
3185 1033
2 14 221 0 0 4224 0 109 119 0 0 4
2893 343
2893 767
3093 767
3093 1033
3 8 222 0 0 4224 0 109 118 0 0 4
2881 343
2881 782
2997 782
2997 1033
1 18 223 0 0 4224 0 109 118 0 0 4
2869 343
2869 787
2907 787
2907 1033
3 2 224 0 0 12416 0 107 108 0 0 5
2935 292
2936 292
2936 288
2921 288
2921 273
5 1 225 0 0 8320 0 109 108 0 0 4
2887 292
2887 288
2903 288
2903 273
3 7 226 0 0 12416 0 55 121 0 0 5
2855 343
2856 343
2856 849
3449 849
3449 1034
2 17 227 0 0 12416 0 55 121 0 0 5
2846 343
2847 343
2847 849
3359 849
3359 1034
1 11 228 0 0 8320 0 55 120 0 0 5
2837 343
2838 343
2838 849
3266 849
3266 1033
4 21 229 0 0 8320 0 110 120 0 0 4
2816 344
2816 687
3176 687
3176 1033
2 15 230 0 0 4224 0 110 119 0 0 4
2804 344
2804 712
3084 712
3084 1033
3 9 231 0 0 4224 0 110 118 0 0 4
2792 344
2792 1015
2988 1015
2988 1033
1 19 232 0 0 4224 0 110 118 0 0 6
2780 344
2780 790
2902 790
2902 1025
2898 1025
2898 1033
5 1 233 0 0 12416 0 110 111 0 0 4
2798 293
2798 289
2809 289
2809 210
3 8 234 0 0 12416 0 56 121 0 0 5
2747 345
2748 345
2748 847
3440 847
3440 1034
2 18 235 0 0 12416 0 56 121 0 0 5
2738 345
2739 345
2739 847
3350 847
3350 1034
1 12 236 0 0 12416 0 56 120 0 0 5
2729 345
2730 345
2730 847
3257 847
3257 1033
4 22 237 0 0 8320 0 112 120 0 0 4
2708 345
2708 690
3167 690
3167 1033
2 16 238 0 0 8320 0 112 119 0 0 4
2696 345
2696 695
3075 695
3075 1033
3 10 239 0 0 4224 0 112 118 0 0 4
2684 345
2684 1020
2979 1020
2979 1033
1 20 240 0 0 4224 0 112 118 0 0 4
2672 345
2672 1025
2889 1025
2889 1033
3 9 241 0 0 8320 0 59 121 0 0 4
2645 345
2645 763
3431 763
3431 1034
2 19 242 0 0 8320 0 59 121 0 0 4
2636 345
2636 773
3341 773
3341 1034
1 13 243 0 0 8320 0 59 120 0 0 4
2627 345
2627 846
3248 846
3248 1033
4 7 244 0 0 8320 0 114 119 0 0 4
2605 345
2605 778
3156 778
3156 1033
2 17 245 0 0 8320 0 114 119 0 0 4
2593 345
2593 699
3066 699
3066 1033
3 11 246 0 0 8320 0 114 118 0 0 4
2581 345
2581 704
2970 704
2970 1033
1 21 247 0 0 4224 0 114 118 0 0 6
2569 345
2569 709
2862 709
2862 859
2880 859
2880 1033
5 1 248 0 0 12416 0 112 113 0 0 4
2690 294
2690 290
2708 290
2708 212
5 1 249 0 0 12416 0 114 115 0 0 4
2587 294
2587 290
2602 290
2602 212
5 1 250 0 0 12416 0 117 116 0 0 4
2460 300
2460 296
2476 296
2476 214
10 0 74 0 0 8320 0 121 0 0 0 4
3422 1034
3422 384
2518 384
2518 350
20 0 75 0 0 8320 0 121 0 0 0 4
3332 1034
3332 379
2509 379
2509 350
14 0 76 0 0 8320 0 120 0 0 0 4
3239 1033
3239 374
2500 374
2500 350
8 4 251 0 0 8320 0 119 117 0 0 4
3147 1033
3147 370
2478 370
2478 351
18 2 252 0 0 4224 0 119 117 0 0 4
3057 1033
3057 365
2466 365
2466 351
12 3 253 0 0 4224 0 118 117 0 0 4
2961 1033
2961 360
2454 360
2454 351
22 1 254 0 0 12416 0 118 117 0 0 6
2871 1033
2871 923
2447 923
2447 360
2442 360
2442 351
14 1 255 0 0 8320 0 124 43 0 0 4
3389 2237
3389 2895
2568 2895
2568 2925
8 2 256 0 0 8320 0 123 43 0 0 4
3296 2236
3296 2900
2559 2900
2559 2925
18 3 257 0 0 4224 0 123 43 0 0 4
3206 2236
3206 2905
2550 2905
2550 2925
12 1 258 0 0 4224 0 125 51 0 0 4
3114 2236
3114 2908
2529 2908
2529 2923
22 2 259 0 0 4224 0 125 51 0 0 4
3024 2236
3024 2913
2520 2913
2520 2923
16 3 260 0 0 4224 0 126 51 0 0 4
2928 2236
2928 2918
2511 2918
2511 2923
0 1 109 0 0 0 0 0 198 350 0 2
1683 2708
1655 2708
5 2 109 0 0 0 0 188 198 0 0 4
1739 2753
1683 2753
1683 2699
1655 2699
4 0 7 0 0 4224 0 129 0 0 0 2
873 2122
601 2122
5 0 4 0 0 4224 0 127 0 0 0 2
871 2009
604 2009
5 0 10 0 0 4224 0 128 0 0 0 2
873 1907
605 1907
4 0 11 0 0 4224 0 130 0 0 0 2
869 1841
610 1841
0 3 261 0 0 4224 0 0 129 366 0 3
1046 1562
1046 2113
925 2113
0 2 262 0 0 4224 0 0 129 365 0 3
1076 1692
1076 2122
924 2122
0 1 263 0 0 4096 0 0 129 358 0 2
1090 2131
925 2131
0 1 263 0 0 4096 0 0 127 367 0 5
1090 2391
1090 2031
962 2031
962 2022
927 2022
4 2 264 0 0 12416 0 175 127 0 0 4
1195 1896
1144 1896
1144 2013
927 2013
0 3 265 0 0 4224 0 0 127 372 0 3
1117 1789
1117 2004
927 2004
0 4 262 0 0 0 0 0 127 369 0 3
1102 1832
1102 1995
927 1995
4 1 266 0 0 8320 0 155 128 0 0 4
1215 2516
982 2516
982 1920
923 1920
2 0 267 0 0 4096 0 128 0 0 370 2
923 1911
946 1911
3 0 265 0 0 0 0 128 0 0 372 3
923 1902
1040 1902
1040 1789
0 2 262 0 0 0 0 0 133 369 0 6
1128 1692
1026 1692
1026 1552
973 1552
973 1562
923 1562
3 4 261 0 0 0 0 136 128 0 0 6
1124 1539
1130 1539
1130 1562
990 1562
990 1893
923 1893
4 1 263 0 0 8320 0 159 130 0 0 4
1210 2391
1030 2391
1030 1850
921 1850
2 0 268 0 0 4096 0 130 0 0 376 2
920 1841
1063 1841
3 3 262 0 0 0 0 130 135 0 0 4
921 1832
1128 1832
1128 1663
1122 1663
4 1 267 0 0 8320 0 163 132 0 0 4
1207 2270
946 2270
946 1655
919 1655
4 2 269 0 0 8320 0 167 132 0 0 4
1203 2143
941 2143
941 1637
919 1637
3 1 265 0 0 0 0 134 131 0 0 4
1127 1789
921 1789
921 1718
913 1718
2 0 12 0 0 4224 0 131 0 0 0 2
877 1718
604 1718
3 0 15 0 0 4224 0 132 0 0 0 2
867 1646
605 1646
3 0 17 0 0 4224 0 133 0 0 0 2
871 1571
594 1571
4 1 268 0 0 8320 0 171 133 0 0 4
1199 2021
1063 2021
1063 1580
923 1580
4 1 270 0 0 16512 0 147 136 0 0 6
1217 2767
1181 2767
1181 2726
1274 2726
1274 1548
1170 1548
4 1 271 0 0 16512 0 143 135 0 0 8
1220 2891
1181 2891
1181 2841
1290 2841
1290 1704
1248 1704
1248 1672
1168 1672
3 1 272 0 0 16512 0 137 134 0 0 8
1218 3015
1183 3015
1183 2968
1310 2968
1310 1833
1219 1833
1219 1798
1173 1798
5 1 273 0 0 4224 0 139 137 0 0 4
1329 3018
1286 3018
1286 3024
1264 3024
4 2 274 0 0 12416 0 179 134 0 0 4
1192 1776
1195 1776
1195 1780
1173 1780
4 2 275 0 0 12416 0 183 135 0 0 4
1191 1650
1190 1650
1190 1654
1168 1654
4 2 276 0 0 12416 0 184 136 0 0 4
1188 1520
1192 1520
1192 1530
1170 1530
0 0 277 0 0 4096 0 0 0 680 702 2
2385 694
2385 719
2 5 278 0 0 4224 0 137 138 0 0 4
1264 3006
1322 3006
1322 2971
1328 2971
1 7 279 0 0 8320 0 139 198 0 0 4
1380 3036
1511 3036
1511 2753
1579 2753
3 8 280 0 0 8320 0 139 198 0 0 4
1380 3024
1556 3024
1556 2744
1579 2744
2 9 281 0 0 8320 0 139 198 0 0 4
1380 3012
1521 3012
1521 2735
1579 2735
4 10 282 0 0 8320 0 139 198 0 0 4
1380 3000
1461 3000
1461 2726
1579 2726
1 11 283 0 0 8320 0 138 198 0 0 4
1379 2989
1486 2989
1486 2717
1579 2717
3 12 284 0 0 8320 0 138 198 0 0 4
1379 2977
1526 2977
1526 2708
1579 2708
2 13 285 0 0 8320 0 138 198 0 0 4
1379 2965
1531 2965
1531 2699
1579 2699
4 14 286 0 0 8320 0 138 198 0 0 4
1379 2953
1466 2953
1466 2690
1579 2690
1 15 287 0 0 8320 0 142 198 0 0 4
1376 2941
1561 2941
1561 2681
1579 2681
2 16 288 0 0 8320 0 142 198 0 0 4
1376 2923
1491 2923
1491 2672
1579 2672
1 17 289 0 0 8320 0 141 198 0 0 4
1374 2911
1541 2911
1541 2663
1579 2663
3 18 290 0 0 8320 0 141 198 0 0 4
1374 2899
1546 2899
1546 2654
1579 2654
2 19 291 0 0 8320 0 141 198 0 0 4
1374 2887
1501 2887
1501 2645
1579 2645
4 20 292 0 0 8320 0 141 198 0 0 4
1374 2875
1536 2875
1536 2636
1579 2636
1 21 293 0 0 8320 0 140 198 0 0 4
1373 2864
1551 2864
1551 2627
1579 2627
3 22 294 0 0 8320 0 140 198 0 0 4
1373 2852
1566 2852
1566 2618
1579 2618
2 7 295 0 0 8320 0 140 199 0 0 4
1373 2840
1470 2840
1470 2590
1578 2590
4 8 296 0 0 8320 0 140 199 0 0 4
1373 2828
1505 2828
1505 2581
1578 2581
1 9 297 0 0 8320 0 146 199 0 0 4
1373 2817
1515 2817
1515 2572
1578 2572
2 10 298 0 0 8320 0 146 199 0 0 4
1373 2799
1475 2799
1475 2563
1578 2563
1 11 299 0 0 8320 0 145 199 0 0 4
1371 2787
1495 2787
1495 2554
1578 2554
3 12 300 0 0 8320 0 145 199 0 0 4
1371 2775
1570 2775
1570 2545
1578 2545
2 13 301 0 0 8320 0 145 199 0 0 4
1371 2763
1480 2763
1480 2536
1578 2536
4 14 302 0 0 8320 0 145 199 0 0 4
1371 2751
1510 2751
1510 2527
1578 2527
1 15 303 0 0 8320 0 144 199 0 0 4
1370 2740
1555 2740
1555 2518
1578 2518
3 16 304 0 0 8320 0 144 199 0 0 4
1370 2728
1520 2728
1520 2509
1578 2509
2 17 305 0 0 8320 0 144 199 0 0 4
1370 2716
1485 2716
1485 2500
1578 2500
4 18 306 0 0 8320 0 144 199 0 0 4
1370 2704
1525 2704
1525 2491
1578 2491
1 19 307 0 0 8320 0 150 199 0 0 4
1373 2692
1530 2692
1530 2482
1578 2482
2 20 308 0 0 8320 0 150 199 0 0 4
1373 2674
1560 2674
1560 2473
1578 2473
1 21 309 0 0 8320 0 149 199 0 0 4
1371 2662
1540 2662
1540 2464
1578 2464
3 22 310 0 0 8320 0 149 199 0 0 4
1371 2650
1545 2650
1545 2455
1578 2455
2 7 311 0 0 8320 0 149 197 0 0 4
1371 2638
1500 2638
1500 2425
1578 2425
4 8 312 0 0 8320 0 149 197 0 0 4
1371 2626
1550 2626
1550 2416
1578 2416
1 9 313 0 0 8320 0 148 197 0 0 4
1370 2615
1565 2615
1565 2407
1578 2407
3 10 314 0 0 8320 0 148 197 0 0 4
1370 2603
1490 2603
1490 2398
1578 2398
2 11 315 0 0 8320 0 148 197 0 0 4
1370 2591
1535 2591
1535 2389
1578 2389
4 12 316 0 0 8320 0 148 197 0 0 4
1370 2579
1505 2579
1505 2380
1578 2380
1 13 317 0 0 8320 0 154 197 0 0 4
1371 2566
1515 2566
1515 2371
1578 2371
2 14 318 0 0 8320 0 154 197 0 0 4
1371 2548
1495 2548
1495 2362
1578 2362
1 15 319 0 0 4224 0 153 197 0 0 4
1369 2536
1570 2536
1570 2353
1578 2353
3 16 320 0 0 8320 0 153 197 0 0 4
1369 2524
1510 2524
1510 2344
1578 2344
2 17 321 0 0 4224 0 153 197 0 0 4
1369 2512
1555 2512
1555 2335
1578 2335
4 18 322 0 0 8320 0 153 197 0 0 4
1369 2500
1520 2500
1520 2326
1578 2326
1 19 323 0 0 8320 0 152 197 0 0 4
1368 2489
1525 2489
1525 2317
1578 2317
3 20 324 0 0 8320 0 152 197 0 0 4
1368 2477
1530 2477
1530 2308
1578 2308
2 21 325 0 0 4224 0 152 197 0 0 4
1368 2465
1560 2465
1560 2299
1578 2299
4 22 326 0 0 4224 0 152 197 0 0 4
1368 2453
1540 2453
1540 2290
1578 2290
1 7 327 0 0 8320 0 158 196 0 0 4
1366 2441
1544 2441
1544 2262
1577 2262
2 8 328 0 0 8320 0 158 196 0 0 4
1366 2423
1499 2423
1499 2253
1577 2253
1 9 329 0 0 4224 0 157 196 0 0 4
1364 2411
1549 2411
1549 2244
1577 2244
3 10 330 0 0 4224 0 157 196 0 0 4
1364 2399
1564 2399
1564 2235
1577 2235
2 11 331 0 0 4224 0 157 196 0 0 4
1364 2387
1534 2387
1534 2226
1577 2226
4 12 332 0 0 8320 0 157 196 0 0 4
1364 2375
1504 2375
1504 2217
1577 2217
1 13 333 0 0 8320 0 156 196 0 0 4
1363 2364
1514 2364
1514 2208
1577 2208
3 14 334 0 0 4224 0 156 196 0 0 4
1363 2352
1569 2352
1569 2199
1577 2199
2 15 335 0 0 8320 0 156 196 0 0 4
1363 2340
1509 2340
1509 2190
1577 2190
4 16 336 0 0 4224 0 156 196 0 0 4
1363 2328
1554 2328
1554 2181
1577 2181
1 17 337 0 0 4224 0 162 196 0 0 4
1363 2320
1519 2320
1519 2172
1577 2172
2 18 338 0 0 4224 0 162 196 0 0 4
1363 2302
1524 2302
1524 2163
1577 2163
1 19 339 0 0 4224 0 161 196 0 0 4
1361 2290
1559 2290
1559 2154
1577 2154
3 20 340 0 0 4224 0 161 196 0 0 4
1361 2278
1539 2278
1539 2145
1577 2145
2 21 341 0 0 4224 0 161 196 0 0 4
1361 2266
1529 2266
1529 2136
1577 2136
4 22 342 0 0 4224 0 161 196 0 0 4
1361 2254
1544 2254
1544 2127
1577 2127
1 7 343 0 0 4224 0 160 201 0 0 4
1360 2243
1550 2243
1550 2094
1578 2094
3 8 344 0 0 4224 0 160 201 0 0 4
1360 2231
1565 2231
1565 2085
1578 2085
2 9 345 0 0 4224 0 160 201 0 0 4
1360 2219
1535 2219
1535 2076
1578 2076
4 10 346 0 0 4224 0 160 201 0 0 4
1360 2207
1515 2207
1515 2067
1578 2067
1 11 347 0 0 4224 0 166 201 0 0 4
1359 2193
1570 2193
1570 2058
1578 2058
2 12 348 0 0 4224 0 166 201 0 0 4
1359 2175
1555 2175
1555 2049
1578 2049
1 13 349 0 0 4224 0 165 201 0 0 4
1357 2163
1520 2163
1520 2040
1578 2040
3 14 350 0 0 4224 0 165 201 0 0 4
1357 2151
1560 2151
1560 2031
1578 2031
2 15 351 0 0 4224 0 165 201 0 0 4
1357 2139
1540 2139
1540 2022
1578 2022
4 16 352 0 0 4224 0 165 201 0 0 4
1357 2127
1530 2127
1530 2013
1578 2013
1 17 353 0 0 4224 0 164 201 0 0 4
1356 2116
1525 2116
1525 2004
1578 2004
3 18 354 0 0 4224 0 164 201 0 0 4
1356 2104
1545 2104
1545 1995
1578 1995
2 19 355 0 0 4224 0 164 201 0 0 4
1356 2092
1550 2092
1550 1986
1578 1986
4 20 356 0 0 4224 0 164 201 0 0 4
1356 2080
1565 2080
1565 1977
1578 1977
1 21 357 0 0 4224 0 170 201 0 0 4
1355 2071
1535 2071
1535 1968
1578 1968
2 22 358 0 0 4224 0 170 201 0 0 4
1355 2053
1570 2053
1570 1959
1578 1959
1 7 359 0 0 4224 0 169 200 0 0 4
1353 2041
1554 2041
1554 1931
1577 1931
3 8 360 0 0 4224 0 169 200 0 0 4
1353 2029
1559 2029
1559 1922
1577 1922
2 9 361 0 0 4224 0 169 200 0 0 4
1353 2017
1539 2017
1539 1913
1577 1913
4 10 362 0 0 4224 0 169 200 0 0 4
1353 2005
1529 2005
1529 1904
1577 1904
1 11 363 0 0 4224 0 168 200 0 0 4
1352 1994
1544 1994
1544 1895
1577 1895
3 12 364 0 0 4224 0 168 200 0 0 4
1352 1982
1549 1982
1549 1886
1577 1886
2 13 365 0 0 4224 0 168 200 0 0 4
1352 1970
1564 1970
1564 1877
1577 1877
4 14 366 0 0 4224 0 168 200 0 0 4
1352 1958
1534 1958
1534 1868
1577 1868
1 15 367 0 0 4224 0 174 200 0 0 4
1351 1946
1569 1946
1569 1859
1577 1859
2 16 368 0 0 4224 0 174 200 0 0 4
1351 1928
1554 1928
1554 1850
1577 1850
1 17 369 0 0 4224 0 173 200 0 0 4
1349 1916
1559 1916
1559 1841
1577 1841
3 18 370 0 0 4224 0 173 200 0 0 4
1349 1904
1539 1904
1539 1832
1577 1832
2 19 371 0 0 4224 0 173 200 0 0 4
1349 1892
1544 1892
1544 1823
1577 1823
4 20 372 0 0 4224 0 173 200 0 0 4
1349 1880
1549 1880
1549 1814
1577 1814
1 21 373 0 0 4224 0 172 200 0 0 4
1348 1869
1564 1869
1564 1805
1577 1805
3 22 374 0 0 4224 0 172 200 0 0 4
1348 1857
1569 1857
1569 1796
1577 1796
2 7 375 0 0 4224 0 172 202 0 0 4
1348 1845
1554 1845
1554 1766
1577 1766
4 8 376 0 0 4224 0 172 202 0 0 4
1348 1833
1559 1833
1559 1757
1577 1757
1 9 377 0 0 4224 0 178 202 0 0 4
1348 1826
1539 1826
1539 1748
1577 1748
2 10 378 0 0 4224 0 178 202 0 0 4
1348 1808
1544 1808
1544 1739
1577 1739
1 11 379 0 0 4224 0 177 202 0 0 4
1346 1796
1564 1796
1564 1730
1577 1730
3 12 380 0 0 4224 0 177 202 0 0 4
1346 1784
1569 1784
1569 1721
1577 1721
2 13 381 0 0 4224 0 177 202 0 0 4
1346 1772
1549 1772
1549 1712
1577 1712
4 14 382 0 0 4224 0 177 202 0 0 4
1346 1760
1554 1760
1554 1703
1577 1703
1 15 383 0 0 4224 0 176 202 0 0 4
1345 1749
1559 1749
1559 1694
1577 1694
16 3 384 0 0 4224 0 202 176 0 0 4
1577 1685
1355 1685
1355 1737
1345 1737
2 17 385 0 0 4224 0 176 202 0 0 4
1345 1725
1564 1725
1564 1676
1577 1676
4 18 386 0 0 4224 0 176 202 0 0 4
1345 1713
1569 1713
1569 1667
1577 1667
1 19 387 0 0 4224 0 182 202 0 0 4
1347 1700
1554 1700
1554 1658
1577 1658
2 20 388 0 0 4224 0 182 202 0 0 4
1347 1682
1559 1682
1559 1649
1577 1649
1 21 389 0 0 4224 0 181 202 0 0 4
1345 1670
1564 1670
1564 1640
1577 1640
3 22 390 0 0 4224 0 181 202 0 0 4
1345 1658
1569 1658
1569 1631
1577 1631
2 7 391 0 0 4224 0 181 203 0 0 4
1345 1646
1558 1646
1558 1603
1576 1603
4 8 392 0 0 4224 0 181 203 0 0 4
1345 1634
1563 1634
1563 1594
1576 1594
1 9 393 0 0 4224 0 180 203 0 0 4
1344 1623
1553 1623
1553 1585
1576 1585
3 10 394 0 0 4224 0 180 203 0 0 4
1344 1611
1568 1611
1568 1576
1576 1576
2 11 395 0 0 4224 0 180 203 0 0 4
1344 1599
1558 1599
1558 1567
1576 1567
4 12 396 0 0 4224 0 180 203 0 0 4
1344 1587
1563 1587
1563 1558
1576 1558
1 13 397 0 0 4224 0 185 203 0 0 4
1344 1570
1568 1570
1568 1549
1576 1549
2 14 398 0 0 4224 0 185 203 0 0 4
1344 1552
1563 1552
1563 1540
1576 1540
1 15 399 0 0 4224 0 186 203 0 0 4
1342 1540
1568 1540
1568 1531
1576 1531
3 16 400 0 0 4224 0 186 203 0 0 4
1342 1528
1568 1528
1568 1522
1576 1522
2 17 401 0 0 4224 0 186 203 0 0 4
1342 1516
1568 1516
1568 1513
1576 1513
4 18 402 0 0 4224 0 186 203 0 0 2
1342 1504
1576 1504
1 19 403 0 0 4224 0 187 203 0 0 4
1341 1493
1568 1493
1568 1495
1576 1495
3 20 404 0 0 4224 0 187 203 0 0 4
1341 1481
1568 1481
1568 1486
1576 1486
21 2 405 0 0 4224 0 203 187 0 0 4
1576 1477
1351 1477
1351 1469
1341 1469
4 22 406 0 0 4224 0 187 203 0 0 4
1341 1457
1568 1457
1568 1468
1576 1468
1 3 407 0 0 4224 0 143 142 0 0 4
1266 2900
1319 2900
1319 2932
1325 2932
5 2 408 0 0 4224 0 141 143 0 0 4
1323 2893
1288 2893
1288 2891
1265 2891
3 5 409 0 0 4224 0 143 140 0 0 4
1266 2882
1316 2882
1316 2846
1322 2846
1 3 410 0 0 4224 0 147 146 0 0 4
1263 2776
1316 2776
1316 2808
1322 2808
5 2 411 0 0 4224 0 145 147 0 0 4
1320 2769
1285 2769
1285 2767
1262 2767
3 5 412 0 0 4224 0 147 144 0 0 4
1263 2758
1313 2758
1313 2722
1319 2722
1 3 413 0 0 4224 0 151 150 0 0 4
1263 2651
1316 2651
1316 2683
1322 2683
5 2 414 0 0 4224 0 149 151 0 0 4
1320 2644
1285 2644
1285 2642
1262 2642
3 5 415 0 0 4224 0 151 148 0 0 4
1263 2633
1313 2633
1313 2597
1319 2597
1 3 416 0 0 4224 0 155 154 0 0 4
1261 2525
1314 2525
1314 2557
1320 2557
5 2 417 0 0 4224 0 153 155 0 0 4
1318 2518
1283 2518
1283 2516
1260 2516
3 5 418 0 0 4224 0 155 152 0 0 4
1261 2507
1311 2507
1311 2471
1317 2471
1 3 419 0 0 4224 0 159 158 0 0 4
1256 2400
1309 2400
1309 2432
1315 2432
5 2 420 0 0 4224 0 157 159 0 0 4
1313 2393
1278 2393
1278 2391
1255 2391
3 5 421 0 0 4224 0 159 156 0 0 4
1256 2382
1306 2382
1306 2346
1312 2346
1 3 422 0 0 4224 0 163 162 0 0 4
1253 2279
1306 2279
1306 2311
1312 2311
5 2 423 0 0 4224 0 161 163 0 0 4
1310 2272
1275 2272
1275 2270
1252 2270
3 5 424 0 0 4224 0 163 160 0 0 4
1253 2261
1303 2261
1303 2225
1309 2225
1 3 425 0 0 4224 0 167 166 0 0 4
1249 2152
1302 2152
1302 2184
1308 2184
5 2 426 0 0 4224 0 165 167 0 0 4
1306 2145
1271 2145
1271 2143
1248 2143
3 5 427 0 0 4224 0 167 164 0 0 4
1249 2134
1299 2134
1299 2098
1305 2098
1 3 428 0 0 4224 0 171 170 0 0 4
1245 2030
1298 2030
1298 2062
1304 2062
5 2 429 0 0 4224 0 169 171 0 0 4
1302 2023
1267 2023
1267 2021
1244 2021
3 5 430 0 0 4224 0 171 168 0 0 4
1245 2012
1295 2012
1295 1976
1301 1976
1 3 431 0 0 4224 0 175 174 0 0 4
1241 1905
1294 1905
1294 1937
1300 1937
5 2 432 0 0 4224 0 173 175 0 0 4
1298 1898
1263 1898
1263 1896
1240 1896
3 5 433 0 0 4224 0 175 172 0 0 4
1241 1887
1291 1887
1291 1851
1297 1851
1 3 434 0 0 4224 0 179 178 0 0 4
1238 1785
1291 1785
1291 1817
1297 1817
5 2 435 0 0 4224 0 177 179 0 0 4
1295 1778
1260 1778
1260 1776
1237 1776
3 5 436 0 0 4224 0 179 176 0 0 4
1238 1767
1288 1767
1288 1731
1294 1731
1 3 437 0 0 4224 0 183 182 0 0 4
1237 1659
1290 1659
1290 1691
1296 1691
5 2 438 0 0 4224 0 181 183 0 0 4
1294 1652
1259 1652
1259 1650
1236 1650
3 5 439 0 0 4224 0 183 180 0 0 4
1237 1641
1287 1641
1287 1605
1293 1605
1 3 440 0 0 4224 0 184 185 0 0 4
1234 1529
1287 1529
1287 1561
1293 1561
5 2 441 0 0 4224 0 186 184 0 0 4
1291 1522
1256 1522
1256 1520
1233 1520
3 5 442 0 0 4224 0 184 187 0 0 4
1234 1511
1284 1511
1284 1475
1290 1475
1 0 443 0 0 4096 0 192 0 0 650 2
1776 2109
2501 2109
2 0 444 0 0 4096 0 192 0 0 669 2
1776 2100
2618 2100
3 0 445 0 0 4096 0 192 0 0 666 2
1776 2091
2753 2091
1 0 446 0 0 4096 0 193 0 0 670 2
1774 1946
2519 1946
2 0 444 0 0 4096 0 193 0 0 669 2
1774 1937
2618 1937
3 0 445 0 0 4096 0 193 0 0 666 2
1774 1928
2753 1928
1 0 443 0 0 4096 0 194 0 0 671 2
1771 1785
2501 1785
2 0 447 0 0 4096 0 194 0 0 668 2
1771 1776
2636 1776
3 0 445 0 0 4096 0 194 0 0 666 2
1771 1767
2753 1767
0 0 448 0 0 4224 0 0 0 739 686 3
2027 527
2876 527
2876 717
0 0 449 0 0 4224 0 0 0 738 690 3
2035 514
2761 514
2761 715
0 0 450 0 0 4224 0 0 0 737 694 3
2048 500
2644 500
2644 717
0 0 451 0 0 4224 0 0 0 736 698 3
2065 487
2534 487
2534 718
1 0 446 0 0 4096 0 195 0 0 670 2
1769 1621
2519 1621
2 0 447 0 0 0 0 195 0 0 668 4
1769 1612
2631 1612
2631 1613
2636 1613
3 0 445 0 0 4096 0 195 0 0 666 2
1769 1603
2753 1603
1 0 452 0 0 4096 0 234 0 0 581 2
2035 795
2035 768
2 0 452 0 0 4096 0 233 0 0 581 2
2080 796
2080 768
1 0 452 0 0 0 0 229 0 0 581 2
2155 793
2155 768
2 0 452 0 0 0 0 230 0 0 581 2
2200 794
2200 768
1 0 452 0 0 0 0 225 0 0 581 2
2263 795
2263 768
2 0 452 0 0 0 0 226 0 0 581 2
2308 796
2308 768
1 0 452 0 0 4096 0 221 0 0 581 2
2373 797
2373 768
2 0 452 0 0 4096 0 222 0 0 581 2
2418 798
2418 768
1 0 452 0 0 0 0 217 0 0 581 2
2480 796
2480 768
2 0 452 0 0 0 0 218 0 0 581 2
2525 797
2525 768
1 0 452 0 0 0 0 213 0 0 581 2
2597 795
2597 768
2 0 452 0 0 0 0 214 0 0 581 2
2642 796
2642 768
1 0 452 0 0 0 0 209 0 0 581 2
2714 793
2714 768
0 2 452 0 0 0 0 0 210 581 0 2
2759 768
2759 794
1 0 452 0 0 0 0 205 0 0 581 2
2828 795
2828 768
0 2 452 0 0 16384 0 0 206 769 0 6
1796 240
1796 539
2002 539
2002 768
2873 768
2873 796
1 0 446 0 0 0 0 191 0 0 649 2
1779 2279
2519 2279
2 0 447 0 0 0 0 191 0 0 668 4
1779 2270
2631 2270
2631 2271
2636 2271
2 0 447 0 0 0 0 190 0 0 668 4
1781 2428
2631 2428
2631 2429
2636 2429
1 0 443 0 0 0 0 190 0 0 650 2
1781 2437
2501 2437
1 0 446 0 0 0 0 189 0 0 649 2
1785 2606
2519 2606
2 0 444 0 0 0 0 189 0 0 669 2
1785 2597
2618 2597
3 0 453 0 0 4096 0 191 0 0 667 2
1779 2261
2735 2261
3 0 453 0 0 0 0 190 0 0 667 4
1781 2419
2730 2419
2730 2420
2735 2420
3 0 453 0 0 0 0 189 0 0 667 4
1785 2588
2730 2588
2730 2589
2735 2589
1 0 443 0 0 0 0 188 0 0 650 4
1789 2766
2496 2766
2496 2767
2501 2767
2 0 444 0 0 0 0 188 0 0 669 2
1789 2757
2618 2757
3 0 453 0 0 0 0 188 0 0 667 2
1789 2748
2735 2748
4 0 3 0 0 0 0 188 0 0 664 2
1789 2739
2867 2739
4 0 3 0 0 0 0 189 0 0 664 2
1785 2579
2867 2579
4 0 3 0 0 0 0 190 0 0 664 2
1781 2410
2867 2410
4 0 3 0 0 0 0 191 0 0 664 2
1779 2252
2867 2252
4 0 3 0 0 0 0 192 0 0 664 2
1776 2082
2867 2082
4 0 3 0 0 0 0 193 0 0 664 2
1774 1919
2867 1919
4 0 3 0 0 0 0 194 0 0 664 2
1771 1758
2867 1758
4 0 3 0 0 0 0 195 0 0 664 2
1769 1594
2867 1594
1 0 110 0 0 0 0 199 0 0 603 2
1654 2545
1737 2545
2 5 110 0 0 0 0 199 189 0 0 4
1654 2536
1737 2536
1737 2593
1735 2593
1 0 111 0 0 0 0 197 0 0 605 2
1654 2380
1733 2380
2 5 111 0 0 0 0 197 190 0 0 4
1654 2371
1733 2371
1733 2424
1731 2424
1 0 112 0 0 0 0 196 0 0 607 2
1653 2217
1731 2217
2 5 112 0 0 0 0 196 191 0 0 4
1653 2208
1731 2208
1731 2266
1729 2266
1 0 113 0 0 0 0 201 0 0 609 2
1654 2049
1728 2049
2 5 113 0 0 0 0 201 192 0 0 4
1654 2040
1728 2040
1728 2096
1726 2096
1 0 114 0 0 0 0 200 0 0 611 2
1653 1886
1726 1886
2 5 114 0 0 0 0 200 193 0 0 4
1653 1877
1726 1877
1726 1933
1724 1933
1 0 115 0 0 0 0 202 0 0 613 2
1653 1721
1681 1721
5 2 115 0 0 0 0 194 202 0 0 4
1721 1772
1681 1772
1681 1712
1653 1712
0 1 116 0 0 0 0 0 203 615 0 3
1680 1608
1680 1558
1652 1558
5 2 116 0 0 0 0 195 203 0 0 4
1719 1608
1680 1608
1680 1549
1652 1549
0 3 119 0 0 0 0 0 198 672 0 4
2412 2704
1678 2704
1678 2672
1649 2672
0 4 79 0 0 0 0 0 198 674 0 4
2302 2713
1673 2713
1673 2663
1649 2663
0 5 118 0 0 0 0 0 198 676 0 4
2194 2722
1668 2722
1668 2654
1649 2654
0 6 117 0 0 0 0 0 198 653 0 4
2074 2731
1663 2731
1663 2645
1649 2645
0 3 119 0 0 0 0 0 199 672 0 4
2412 2541
1677 2541
1677 2509
1648 2509
0 4 79 0 0 0 0 0 199 674 0 4
2302 2550
1672 2550
1672 2500
1648 2500
0 5 118 0 0 0 0 0 199 676 0 4
2194 2559
1667 2559
1667 2491
1648 2491
0 6 117 0 0 0 0 0 199 653 0 4
2074 2568
1662 2568
1662 2482
1648 2482
0 3 119 0 0 0 0 0 197 672 0 4
2412 2376
1677 2376
1677 2344
1648 2344
0 4 79 0 0 0 0 0 197 674 0 4
2302 2385
1672 2385
1672 2335
1648 2335
0 5 118 0 0 0 0 0 197 676 0 4
2194 2394
1667 2394
1667 2326
1648 2326
0 6 117 0 0 0 0 0 197 653 0 4
2074 2403
1662 2403
1662 2317
1648 2317
0 3 119 0 0 0 0 0 196 672 0 4
2412 2213
1676 2213
1676 2181
1647 2181
0 4 79 0 0 0 0 0 196 674 0 4
2302 2222
1671 2222
1671 2172
1647 2172
0 5 118 0 0 0 0 0 196 676 0 4
2194 2231
1666 2231
1666 2163
1647 2163
0 6 117 0 0 0 0 0 196 653 0 4
2074 2240
1661 2240
1661 2154
1647 2154
0 3 119 0 0 0 0 0 201 672 0 4
2412 2045
1677 2045
1677 2013
1648 2013
0 4 79 0 0 0 0 0 201 674 0 4
2302 2054
1672 2054
1672 2004
1648 2004
0 5 118 0 0 0 0 0 201 676 0 4
2194 2063
1667 2063
1667 1995
1648 1995
0 6 117 0 0 0 0 0 201 653 0 4
2074 2072
1662 2072
1662 1986
1648 1986
0 3 119 0 0 0 0 0 200 672 0 4
2412 1882
1676 1882
1676 1850
1647 1850
0 4 79 0 0 0 0 0 200 674 0 4
2302 1891
1671 1891
1671 1841
1647 1841
0 5 118 0 0 0 0 0 200 676 0 4
2194 1900
1666 1900
1666 1832
1647 1832
0 6 117 0 0 0 0 0 200 678 0 4
2074 1909
1661 1909
1661 1823
1647 1823
0 3 119 0 0 0 0 0 202 672 0 4
2412 1717
1676 1717
1676 1685
1647 1685
0 4 79 0 0 0 0 0 202 674 0 4
2302 1726
1671 1726
1671 1676
1647 1676
0 5 118 0 0 0 0 0 202 676 0 4
2194 1735
1666 1735
1666 1667
1647 1667
0 6 117 0 0 0 0 0 202 678 0 4
2074 1744
1661 1744
1661 1658
1647 1658
0 3 119 0 0 0 0 0 203 672 0 4
2412 1554
1675 1554
1675 1522
1646 1522
0 4 79 0 0 0 0 0 203 674 0 4
2302 1563
1670 1563
1670 1513
1646 1513
0 5 118 0 0 0 0 0 203 676 0 4
2194 1572
1665 1572
1665 1504
1646 1504
0 6 117 0 0 0 0 0 203 678 0 4
2074 1582
1660 1582
1660 1495
1646 1495
0 0 454 0 0 4224 0 0 0 654 0 2
2849 1979
2849 2787
0 0 446 0 0 4096 0 0 0 670 0 2
2519 1981
2519 2791
0 0 443 0 0 4096 0 0 0 671 0 2
2501 1984
2501 2786
0 0 455 0 0 4224 0 0 0 655 0 2
2284 1979
2284 2784
0 0 456 0 0 4224 0 0 0 656 0 2
2176 1976
2176 2786
0 0 117 0 0 0 0 0 0 678 0 2
2074 1983
2074 2783
0 0 454 0 0 0 0 0 0 665 0 2
2849 1697
2849 1983
0 0 455 0 0 0 0 0 0 675 0 2
2284 1707
2284 1984
0 0 456 0 0 0 0 0 0 677 0 2
2176 1697
2176 1980
7 0 27 0 0 20608 0 244 0 0 0 6
677 245
677 281
765 281
765 1040
775 1040
775 2228
6 0 28 0 0 20608 0 244 0 0 0 6
671 245
671 289
755 289
755 1047
765 1047
765 2229
5 0 29 0 0 20608 0 244 0 0 0 6
665 245
665 295
746 295
746 1054
755 1054
755 2230
4 0 30 0 0 20608 0 244 0 0 0 6
659 245
659 303
735 303
735 1056
745 1056
745 2230
3 0 31 0 0 28800 0 244 0 0 0 8
653 245
653 325
685 325
685 412
725 412
725 1063
735 1063
735 2232
2 0 32 0 0 20608 0 244 0 0 0 6
647 245
647 356
702 356
702 1071
725 1071
725 2230
1 0 33 0 0 12416 0 244 0 0 0 4
641 245
641 405
792 405
792 2231
4 0 3 0 0 4224 0 204 0 0 0 2
2867 912
2867 2781
3 0 454 0 0 0 0 204 0 0 0 2
2849 918
2849 1703
4 0 445 0 0 4224 0 208 0 0 0 2
2753 910
2753 2787
3 0 453 0 0 4224 0 208 0 0 0 2
2735 916
2735 2787
4 0 447 0 0 4224 0 212 0 0 0 2
2636 912
2636 2810
3 0 444 0 0 4224 0 212 0 0 0 2
2618 918
2618 2799
4 0 446 0 0 4224 0 216 0 0 0 2
2519 913
2519 1987
3 0 443 0 0 4224 0 216 0 0 0 2
2501 919
2501 1989
4 0 119 0 0 4224 0 220 0 0 0 2
2412 914
2412 2786
3 0 457 0 0 4224 0 220 0 0 0 2
2394 920
2394 2789
4 0 79 0 0 4224 0 224 0 0 0 2
2302 912
2302 2786
3 0 455 0 0 0 0 224 0 0 0 2
2284 918
2284 1713
4 0 118 0 0 4224 0 228 0 0 0 2
2194 910
2194 2781
3 0 456 0 0 0 0 228 0 0 0 2
2176 916
2176 1702
4 0 117 0 0 4224 0 235 0 0 0 2
2074 912
2074 1987
3 0 458 0 0 4224 0 235 0 0 0 2
2056 918
2056 2786
0 0 277 0 0 8320 0 0 0 744 0 4
1951 261
1951 694
2419 694
2419 720
0 0 459 0 0 4224 0 0 0 743 706 4
1958 270
1958 677
2306 677
2306 717
0 0 460 0 0 4224 0 0 0 742 710 4
1970 279
1970 665
2207 665
2207 715
0 0 461 0 0 4096 0 0 0 741 714 4
1979 288
1979 658
2090 658
2090 717
3 2 462 0 0 8320 0 205 204 0 0 4
2819 840
2819 855
2849 855
2849 864
3 1 463 0 0 8320 0 206 204 0 0 4
2882 841
2882 855
2867 855
2867 864
1 1 448 0 0 0 0 207 206 0 0 4
2812 721
2812 717
2891 717
2891 796
2 2 464 0 0 4224 0 207 205 0 0 4
2812 757
2812 787
2810 787
2810 795
3 2 465 0 0 8320 0 209 208 0 0 4
2705 838
2705 853
2735 853
2735 862
3 1 466 0 0 8320 0 210 208 0 0 4
2768 839
2768 853
2753 853
2753 862
1 1 449 0 0 0 0 211 210 0 0 4
2698 719
2698 715
2777 715
2777 794
2 2 467 0 0 4224 0 211 209 0 0 4
2698 755
2698 785
2696 785
2696 793
3 2 468 0 0 8320 0 213 212 0 0 4
2588 840
2588 855
2618 855
2618 864
3 1 469 0 0 8320 0 214 212 0 0 4
2651 841
2651 855
2636 855
2636 864
1 1 450 0 0 0 0 215 214 0 0 4
2581 721
2581 717
2660 717
2660 796
2 2 470 0 0 4224 0 215 213 0 0 4
2581 757
2581 787
2579 787
2579 795
3 2 471 0 0 8320 0 217 216 0 0 4
2471 841
2471 856
2501 856
2501 865
3 1 472 0 0 8320 0 218 216 0 0 4
2534 842
2534 856
2519 856
2519 865
1 1 451 0 0 0 0 219 218 0 0 4
2464 722
2464 718
2543 718
2543 797
2 2 473 0 0 4224 0 219 217 0 0 4
2464 758
2464 788
2462 788
2462 796
3 2 474 0 0 8320 0 221 220 0 0 4
2364 842
2364 857
2394 857
2394 866
3 1 475 0 0 8320 0 222 220 0 0 4
2427 843
2427 857
2412 857
2412 866
1 1 277 0 0 0 0 223 222 0 0 4
2357 723
2357 719
2436 719
2436 798
2 2 476 0 0 4224 0 223 221 0 0 4
2357 759
2357 789
2355 789
2355 797
3 2 477 0 0 8320 0 225 224 0 0 4
2254 840
2254 855
2284 855
2284 864
3 1 478 0 0 8320 0 226 224 0 0 4
2317 841
2317 855
2302 855
2302 864
1 1 459 0 0 0 0 227 226 0 0 4
2247 721
2247 717
2326 717
2326 796
2 2 479 0 0 4224 0 227 225 0 0 4
2247 757
2247 787
2245 787
2245 795
3 2 480 0 0 8320 0 229 228 0 0 4
2146 838
2146 853
2176 853
2176 862
3 1 481 0 0 8320 0 230 228 0 0 4
2209 839
2209 853
2194 853
2194 862
1 1 460 0 0 0 0 231 230 0 0 4
2139 719
2139 715
2218 715
2218 794
2 2 482 0 0 4224 0 231 229 0 0 4
2139 755
2139 785
2137 785
2137 793
3 2 483 0 0 8320 0 234 235 0 0 4
2026 840
2026 855
2056 855
2056 864
3 1 484 0 0 8320 0 233 235 0 0 4
2089 841
2089 855
2074 855
2074 864
1 1 461 0 0 0 0 232 233 0 0 4
2019 721
2019 717
2098 717
2098 796
2 2 485 0 0 4224 0 232 234 0 0 4
2019 757
2019 787
2017 787
2017 795
4 0 486 0 0 8192 0 239 0 0 724 3
1797 146
1765 146
1765 185
3 2 487 0 0 8320 0 238 239 0 0 4
1875 127
1858 127
1858 164
1845 164
3 1 488 0 0 4224 0 237 239 0 0 4
1873 165
1853 165
1853 146
1845 146
1 0 489 0 0 4096 0 237 0 0 720 2
1918 174
2011 174
1 0 489 0 0 0 0 236 0 0 735 3
1989 133
2011 133
2011 185
2 1 490 0 0 4224 0 236 238 0 0 4
1953 133
1930 133
1930 136
1920 136
0 2 452 0 0 0 0 0 237 723 0 3
1935 157
1935 156
1918 156
0 2 452 0 0 0 0 0 238 769 0 6
1847 240
1914 240
1914 193
1935 193
1935 118
1920 118
0 6 486 0 0 4224 0 0 246 0 0 11
1964 185
1482 185
1482 231
1010 231
1010 282
1011 282
1011 299
836 299
836 312
550 312
550 248
7 0 8 0 0 20608 0 245 0 0 0 6
617 247
617 437
700 437
700 824
453 824
453 2244
6 0 5 0 0 20608 0 245 0 0 0 6
611 247
611 430
687 430
687 816
440 816
440 2241
5 0 9 0 0 20608 0 245 0 0 0 6
605 247
605 423
683 423
683 804
433 804
433 2237
4 0 14 0 0 20608 0 245 0 0 0 6
599 247
599 409
671 409
671 797
423 797
423 2239
3 0 13 0 0 12416 0 245 0 0 0 4
593 247
593 369
411 369
411 2237
2 0 16 0 0 12416 0 245 0 0 0 4
587 247
587 364
406 364
406 2236
1 0 18 0 0 12416 0 245 0 0 0 4
581 247
581 357
399 357
399 2239
1 0 486 0 0 0 0 246 0 0 724 3
520 248
520 290
550 290
5 0 486 0 0 0 0 246 0 0 724 3
544 248
544 274
550 274
4 0 486 0 0 0 0 246 0 0 724 3
538 248
538 285
550 285
14 0 489 0 0 12416 0 240 0 0 0 4
2143 382
2189 382
2189 185
1968 185
0 8 451 0 0 0 0 0 240 838 0 6
1632 622
2065 622
2065 475
2058 475
2058 409
2079 409
0 7 450 0 0 0 0 0 240 839 0 4
1671 607
2048 607
2048 400
2079 400
0 6 449 0 0 0 0 0 240 840 0 4
1708 587
2035 587
2035 391
2079 391
0 5 448 0 0 0 0 0 240 841 0 4
1748 573
2027 573
2027 382
2079 382
10 0 491 0 0 4096 0 241 0 0 758 2
1990 315
1929 315
0 8 461 0 0 0 0 0 241 834 0 6
1446 458
1553 458
1553 408
1890 408
1890 288
1990 288
0 7 460 0 0 0 0 0 241 835 0 6
1457 443
1558 443
1558 415
1882 415
1882 279
1990 279
0 6 459 0 0 0 0 0 241 836 0 4
1470 432
1873 432
1873 270
1990 270
0 5 277 0 0 0 0 0 241 837 0 4
1483 424
1866 424
1866 261
1990 261
1 0 2 0 0 4096 0 240 0 0 757 2
2079 346
1945 346
2 0 491 0 0 4096 0 240 0 0 758 2
2079 355
1929 355
3 0 491 0 0 0 0 240 0 0 758 2
2079 364
1929 364
4 0 2 0 0 0 0 240 0 0 757 2
2079 373
1945 373
11 12 492 0 0 8320 0 240 241 0 0 4
2079 445
2062 445
2062 279
2054 279
13 10 493 0 0 8320 0 241 240 0 0 4
2054 270
2066 270
2066 436
2079 436
14 9 494 0 0 8320 0 241 240 0 0 4
2054 261
2071 261
2071 427
2079 427
4 0 2 0 0 0 0 241 0 0 757 2
1990 252
1945 252
3 0 2 0 0 0 0 241 0 0 757 2
1990 243
1945 243
1 0 2 0 0 0 0 241 0 0 757 2
1990 225
1945 225
2 0 491 0 0 0 0 241 0 0 758 2
1990 234
1929 234
0 0 2 0 0 4224 0 0 0 757 0 2
1945 395
1945 2784
0 0 2 0 0 0 0 0 0 868 0 6
1548 449
1548 433
1633 433
1633 395
1945 395
1945 201
0 0 491 0 0 8320 0 0 0 833 0 3
1326 202
1929 202
1929 2783
10 0 491 0 0 0 0 290 0 0 833 2
1344 180
1326 180
18 10 495 0 0 8320 0 290 288 0 0 4
1408 180
1420 180
1420 400
1488 400
9 0 2 0 0 0 0 246 0 0 763 3
541 170
541 162
571 162
9 0 2 0 0 0 0 245 0 0 763 2
602 169
602 162
0 9 2 0 0 0 0 0 244 764 0 5
556 271
571 271
571 162
662 162
662 167
7 0 2 0 0 0 0 246 0 0 950 7
556 248
556 406
456 406
456 413
446 413
446 408
34 408
3 0 491 0 0 0 0 246 0 0 766 2
532 248
532 259
2 0 491 0 0 0 0 246 0 0 767 3
526 248
526 259
562 259
8 0 491 0 0 0 0 246 0 0 951 5
562 248
562 410
451 410
451 405
13 405
4 1 496 0 0 8320 0 285 243 0 0 4
1831 324
1831 254
743 254
743 231
1 3 452 0 0 8320 0 242 285 0 0 4
769 229
769 240
1849 240
1849 318
1 0 497 0 0 8192 0 247 0 0 901 3
528 15
519 15
519 83
2 0 498 0 0 8320 0 247 0 0 858 3
558 15
563 15
563 83
0 2 497 0 0 8320 0 0 285 792 0 5
1289 1411
1811 1411
1811 444
1849 444
1849 372
3 1 499 0 0 8320 0 249 258 0 0 5
1018 1427
560 1427
560 416
643 416
643 435
3 1 500 0 0 8320 0 250 259 0 0 5
1013 1380
532 1380
532 426
580 426
580 432
3 1 501 0 0 16512 0 251 282 0 0 6
1013 1336
384 1336
384 1055
395 1055
395 417
506 417
3 1 502 0 0 4224 0 252 283 0 0 7
1013 1293
375 1293
375 1048
384 1048
384 410
443 410
443 417
3 1 503 0 0 8320 0 253 279 0 0 7
1013 1251
719 1251
719 317
471 317
471 157
400 157
400 167
3 1 504 0 0 8320 0 254 281 0 0 7
1013 1212
677 1212
677 329
459 329
459 141
326 141
326 147
3 1 505 0 0 8320 0 255 280 0 0 7
1013 1170
693 1170
693 350
442 350
442 127
258 127
258 150
3 1 506 0 0 8320 0 248 278 0 0 7
1015 1129
706 1129
706 341
448 341
448 117
202 117
202 170
1 0 497 0 0 0 0 250 0 0 792 2
1058 1389
1289 1389
1 0 497 0 0 0 0 251 0 0 792 2
1058 1345
1289 1345
1 0 497 0 0 0 0 252 0 0 792 2
1058 1302
1289 1302
1 0 497 0 0 0 0 253 0 0 792 2
1058 1260
1289 1260
1 0 497 0 0 0 0 254 0 0 792 2
1058 1221
1289 1221
2 0 497 0 0 0 0 255 0 0 792 2
1058 1161
1289 1161
1 0 497 0 0 0 0 248 0 0 792 2
1060 1138
1289 1138
0 2 507 0 0 4096 0 0 249 803 0 3
1232 1142
1232 1418
1063 1418
0 2 508 0 0 8192 0 0 251 805 0 4
1224 1112
1204 1112
1204 1327
1058 1327
0 2 509 0 0 8192 0 0 254 808 0 4
1221 1058
1119 1058
1119 1203
1058 1203
0 2 510 0 0 4096 0 0 248 810 0 4
1217 1022
1069 1022
1069 1120
1060 1120
0 1 497 0 0 0 0 0 249 899 0 6
249 462
375 462
375 976
1289 976
1289 1436
1063 1436
2 5 511 0 0 4224 0 256 297 0 0 4
793 731
963 731
963 727
976 727
3 1 512 0 0 8320 0 263 256 0 0 3
639 608
639 731
763 731
2 6 513 0 0 4224 0 257 297 0 0 4
618 710
968 710
968 736
976 736
3 1 514 0 0 4224 0 261 257 0 0 3
576 606
576 710
588 710
1 0 515 0 0 4096 0 262 0 0 798 3
659 513
659 492
643 492
2 2 515 0 0 4224 0 258 263 0 0 4
643 465
643 555
630 555
630 563
2 1 516 0 0 8320 0 262 263 0 0 4
659 549
659 555
648 555
648 563
1 0 517 0 0 4096 0 260 0 0 801 3
596 511
596 490
580 490
2 2 517 0 0 4224 0 259 261 0 0 4
580 462
580 553
567 553
567 561
2 1 518 0 0 8320 0 260 261 0 0 4
596 547
596 553
585 553
585 561
10 0 507 0 0 8320 0 268 0 0 0 3
1622 993
1622 1142
1225 1142
11 2 519 0 0 8320 0 268 250 0 0 5
1631 993
1631 1129
1214 1129
1214 1371
1058 1371
12 0 508 0 0 8320 0 268 0 0 0 3
1640 993
1640 1112
1219 1112
13 2 520 0 0 8320 0 268 252 0 0 5
1649 993
1649 1094
1183 1094
1183 1284
1058 1284
2 2 521 0 0 8320 0 267 253 0 0 5
1465 992
1465 1077
1152 1077
1152 1242
1058 1242
2 0 509 0 0 8320 0 266 0 0 0 3
1489 993
1489 1058
1217 1058
2 1 522 0 0 8320 0 265 255 0 0 5
1515 991
1515 1041
1089 1041
1089 1179
1058 1179
2 0 510 0 0 8320 0 264 0 0 0 3
1542 992
1542 1022
1214 1022
13 1 523 0 0 4224 0 269 264 0 0 4
1523 863
1523 954
1542 954
1542 962
12 1 524 0 0 4224 0 269 265 0 0 4
1514 863
1514 953
1515 953
1515 961
11 1 525 0 0 4224 0 269 266 0 0 4
1505 863
1505 950
1489 950
1489 963
10 1 526 0 0 4224 0 269 267 0 0 4
1496 863
1496 954
1465 954
1465 962
2 8 527 0 0 4224 0 270 268 0 0 4
1632 697
1632 901
1658 901
1658 929
2 7 528 0 0 4224 0 271 268 0 0 4
1671 696
1671 906
1649 906
1649 929
2 6 529 0 0 4224 0 272 268 0 0 4
1708 692
1708 911
1640 911
1640 929
2 5 530 0 0 4224 0 273 268 0 0 4
1748 694
1748 916
1631 916
1631 929
14 9 531 0 0 8320 0 269 268 0 0 4
1550 863
1550 921
1676 921
1676 929
1 0 2 0 0 0 0 269 0 0 823 2
1469 799
1469 785
2 0 2 0 0 0 0 269 0 0 823 2
1478 799
1478 785
3 0 2 0 0 0 0 269 0 0 823 2
1487 799
1487 785
4 0 2 0 0 0 0 269 0 0 827 4
1496 799
1496 785
1428 785
1428 799
1 0 2 0 0 0 0 268 0 0 827 2
1595 929
1595 918
2 0 2 0 0 0 0 268 0 0 827 2
1604 929
1604 918
3 0 2 0 0 0 0 268 0 0 827 2
1613 929
1613 918
0 4 2 0 0 0 0 0 268 950 0 7
34 771
806 771
806 799
1438 799
1438 918
1622 918
1622 929
2 8 532 0 0 4224 0 277 269 0 0 4
1470 694
1470 791
1532 791
1532 799
2 7 533 0 0 12416 0 276 269 0 0 4
1510 696
1510 744
1523 744
1523 799
2 6 534 0 0 12416 0 274 269 0 0 4
1547 692
1547 727
1514 727
1514 799
2 5 535 0 0 8320 0 275 269 0 0 4
1587 694
1587 773
1505 773
1505 799
0 9 491 0 0 0 0 0 269 833 0 3
1446 755
1550 755
1550 799
0 0 491 0 0 0 0 0 0 889 0 6
1326 99
1326 428
1439 428
1439 730
1446 730
1446 762
0 1 461 0 0 0 0 0 277 883 0 3
1446 373
1446 658
1470 658
0 1 460 0 0 0 0 0 276 882 0 4
1457 364
1457 646
1510 646
1510 660
0 1 459 0 0 0 0 0 274 881 0 4
1470 355
1470 639
1547 639
1547 656
0 1 277 0 0 0 0 0 275 880 0 5
1483 346
1483 629
1590 629
1590 658
1587 658
0 1 451 0 0 0 0 0 270 876 0 4
1590 512
1590 622
1632 622
1632 661
0 1 450 0 0 0 0 0 271 875 0 4
1603 503
1603 607
1671 607
1671 660
0 1 449 0 0 0 0 0 272 874 0 4
1615 494
1615 587
1708 587
1708 656
0 1 448 0 0 0 0 0 273 861 0 4
1625 485
1625 573
1748 573
1748 658
2 0 536 0 0 4096 0 279 0 0 937 2
391 168
391 75
2 0 537 0 0 4096 0 280 0 0 938 2
249 151
249 93
2 0 536 0 0 4096 0 278 0 0 937 2
193 170
193 75
3 0 538 0 0 4096 0 278 0 0 935 2
184 170
184 43
4 0 539 0 0 4096 0 278 0 0 934 2
175 170
175 34
5 0 540 0 0 4096 0 278 0 0 922 2
189 220
188 220
3 0 541 0 0 4096 0 279 0 0 936 2
382 167
382 52
3 0 541 0 0 0 0 280 0 0 936 2
240 150
240 52
2 0 538 0 0 0 0 281 0 0 935 4
308 147
308 49
309 49
309 44
4 0 542 0 0 0 0 279 0 0 973 2
391 213
391 213
4 0 543 0 0 0 0 280 0 0 921 2
249 196
249 196
3 0 544 0 0 0 0 281 0 0 976 2
317 193
317 193
2 0 537 0 0 4096 0 282 0 0 938 2
488 417
488 93
3 0 536 0 0 4224 0 283 0 0 937 2
425 417
425 75
2 0 537 0 0 4096 0 283 0 0 938 2
434 418
434 93
4 0 545 0 0 0 0 283 0 0 932 2
434 463
434 463
0 2 498 0 0 0 0 0 291 0 0 2
545 83
571 83
0 0 2 0 0 0 0 0 0 860 950 3
861 480
861 659
34 659
0 0 2 0 0 0 0 0 0 868 867 2
1394 480
802 480
0 5 448 0 0 0 0 0 287 862 0 3
1386 627
1386 485
1635 485
4 1 448 0 0 0 0 284 297 0 0 6
1275 627
1389 627
1389 941
849 941
849 691
976 691
2 0 546 0 0 4096 0 284 0 0 905 2
1227 645
1214 645
10 1 547 0 0 12416 0 297 284 0 0 4
1040 718
1044 718
1044 627
1227 627
12 1 548 0 0 8320 0 287 286 0 0 4
1699 503
1740 503
1740 461
1748 461
0 1 549 0 0 4096 0 0 285 869 0 3
1794 401
1831 401
1831 372
9 0 2 0 0 0 0 326 0 0 0 3
837 420
802 420
802 485
1 0 2 0 0 0 0 287 0 0 0 3
1635 449
1394 449
1394 485
3 0 549 0 0 4224 0 286 0 0 0 2
1794 470
1794 356
13 2 550 0 0 4224 0 287 286 0 0 4
1699 494
1735 494
1735 479
1748 479
14 9 551 0 0 8320 0 288 287 0 0 4
1552 346
1567 346
1567 530
1635 530
13 10 552 0 0 8320 0 288 287 0 0 4
1552 355
1576 355
1576 539
1635 539
12 11 553 0 0 8320 0 288 287 0 0 4
1552 364
1585 364
1585 548
1635 548
6 0 449 0 0 0 0 287 0 0 907 4
1635 494
1395 494
1395 769
1379 769
7 0 450 0 0 0 0 287 0 0 908 4
1635 503
1407 503
1407 782
1350 782
8 0 451 0 0 0 0 287 0 0 909 4
1635 512
1420 512
1420 796
1327 796
11 2 554 0 0 8320 0 290 287 0 0 4
1408 117
1624 117
1624 458
1635 458
12 3 555 0 0 8320 0 290 287 0 0 4
1408 126
1611 126
1611 467
1635 467
13 4 556 0 0 8320 0 290 287 0 0 4
1408 135
1601 135
1601 476
1635 476
5 0 277 0 0 0 0 288 0 0 955 2
1488 346
1149 346
6 0 459 0 0 0 0 288 0 0 956 2
1488 355
1134 355
7 0 460 0 0 0 0 288 0 0 957 2
1488 364
1119 364
8 0 461 0 0 4224 0 288 0 0 958 3
1488 373
1094 373
1094 404
14 1 557 0 0 8320 0 290 288 0 0 4
1408 144
1462 144
1462 310
1488 310
15 2 558 0 0 8320 0 290 288 0 0 4
1408 153
1454 153
1454 319
1488 319
16 3 559 0 0 8320 0 290 288 0 0 4
1408 162
1445 162
1445 328
1488 328
17 4 560 0 0 8320 0 290 288 0 0 4
1408 171
1437 171
1437 337
1488 337
2 0 561 0 0 4224 0 290 0 0 939 2
1344 108
795 108
1 0 491 0 0 0 0 290 0 0 951 4
1338 99
532 99
532 107
13 107
1 9 562 0 0 8320 0 7 290 0 0 3
1048 62
1048 171
1344 171
1 8 563 0 0 8320 0 6 290 0 0 3
1084 61
1084 162
1344 162
1 7 564 0 0 8320 0 1 290 0 0 3
1118 62
1118 153
1344 153
1 6 565 0 0 8320 0 2 290 0 0 3
1151 58
1151 144
1344 144
1 5 566 0 0 8320 0 5 290 0 0 3
1186 60
1186 135
1344 135
1 4 567 0 0 8320 0 3 290 0 0 3
1224 62
1224 126
1344 126
1 3 568 0 0 8320 0 4 290 0 0 3
1264 63
1264 117
1344 117
2 0 491 0 0 0 0 289 0 0 951 2
48 280
13 280
1 0 497 0 0 0 0 289 0 0 901 2
82 280
82 282
0 2 497 0 0 0 0 0 327 901 0 4
144 282
144 440
249 440
249 493
1 0 2 0 0 0 0 327 0 0 950 3
249 529
249 635
34 635
0 0 497 0 0 0 0 0 0 0 0 4
79 282
144 282
144 83
541 83
1 0 541 0 0 0 0 308 0 0 936 4
83 139
106 139
106 140
119 140
2 0 546 0 0 0 0 295 0 0 905 2
1228 734
1215 734
2 0 546 0 0 0 0 296 0 0 905 2
1228 692
1215 692
2 2 546 0 0 4224 0 292 294 0 0 6
1072 611
1214 611
1214 689
1215 689
1215 774
1228 774
0 1 569 0 0 4224 0 0 292 954 0 3
942 169
942 611
1042 611
4 2 449 0 0 0 0 296 297 0 0 6
1276 674
1379 674
1379 920
865 920
865 700
976 700
4 3 450 0 0 0 0 295 297 0 0 6
1276 716
1350 716
1350 889
891 889
891 709
976 709
4 4 451 0 0 0 0 294 297 0 0 6
1276 756
1327 756
1327 860
910 860
910 718
976 718
1 11 570 0 0 4224 0 296 297 0 0 4
1228 674
1053 674
1053 727
1040 727
1 12 571 0 0 4224 0 295 297 0 0 4
1228 716
1048 716
1048 736
1040 736
13 1 572 0 0 4224 0 297 294 0 0 4
1040 745
1220 745
1220 756
1228 756
2 7 573 0 0 12416 0 299 297 0 0 4
567 643
722 643
722 745
976 745
2 8 574 0 0 12416 0 298 297 0 0 4
568 683
680 683
680 754
976 754
14 9 575 0 0 8320 0 326 297 0 0 4
901 420
927 420
927 772
976 772
1 3 576 0 0 4224 0 298 302 0 0 3
538 683
430 683
430 606
3 1 577 0 0 8320 0 300 299 0 0 3
493 608
493 643
537 643
0 0 545 0 0 4096 0 0 0 932 0 3
434 467
456 467
456 455
1 4 578 0 0 4224 0 304 305 0 0 4
669 57
626 57
626 44
618 44
4 2 579 0 0 4224 0 291 304 0 0 4
616 83
661 83
661 75
669 75
0 0 543 0 0 8192 0 0 0 979 0 3
245 223
249 223
249 193
0 0 540 0 0 4096 0 0 0 0 952 3
188 215
188 232
190 232
0 2 537 0 0 0 0 0 328 938 0 4
136 234
136 448
210 448
210 493
0 2 536 0 0 0 0 0 329 937 0 4
127 187
127 459
178 459
178 495
0 2 541 0 0 4224 0 0 330 936 0 4
117 140
117 470
147 470
147 494
0 2 538 0 0 4224 0 0 331 935 0 4
108 100
108 477
116 477
116 494
1 2 539 0 0 4224 0 310 332 0 0 4
90 52
90 475
80 475
80 493
1 0 580 0 0 4096 0 301 0 0 929 3
513 513
513 492
497 492
3 2 580 0 0 4224 0 282 300 0 0 4
497 463
497 555
484 555
484 563
2 1 581 0 0 8320 0 301 300 0 0 4
513 549
513 555
502 555
502 563
1 0 545 0 0 0 0 303 0 0 932 3
450 511
450 490
434 490
3 2 545 0 0 4224 0 0 302 0 0 4
434 460
434 553
421 553
421 561
2 1 582 0 0 8320 0 303 302 0 0 4
450 547
450 553
439 553
439 561
1 1 539 0 0 0 0 310 305 0 0 5
90 52
90 34
179 34
179 35
572 35
1 2 538 0 0 0 0 309 305 0 0 8
85 99
108 99
108 100
108 100
108 43
304 43
304 44
573 44
0 3 541 0 0 0 0 0 305 0 0 6
97 140
119 140
119 52
400 52
400 53
572 53
1 1 536 0 0 0 0 307 291 0 0 6
79 187
127 187
127 75
447 75
447 74
570 74
1 3 537 0 0 12416 0 306 291 0 0 6
80 234
136 234
136 93
505 93
505 92
570 92
3 1 561 0 0 0 0 304 317 0 0 4
715 66
795 66
795 169
803 169
1 0 2 0 0 0 0 332 0 0 950 3
80 529
80 549
34 549
1 0 2 0 0 0 0 331 0 0 950 3
116 530
116 566
34 566
1 0 2 0 0 0 0 330 0 0 950 3
147 530
147 582
34 582
1 0 2 0 0 0 0 329 0 0 950 3
178 531
178 602
34 602
1 0 2 0 0 0 0 328 0 0 950 3
210 529
210 618
34 618
2 0 491 0 0 0 0 310 0 0 951 4
56 52
18 52
18 53
13 53
2 0 491 0 0 0 0 309 0 0 951 4
51 99
28 99
28 100
13 100
2 0 491 0 0 0 0 308 0 0 951 4
49 139
18 139
18 146
13 146
2 0 491 0 0 0 0 307 0 0 951 4
45 187
18 187
18 188
13 188
2 0 491 0 0 0 0 306 0 0 951 2
46 234
13 234
1 0 2 0 0 0 0 311 0 0 0 2
34 781
34 11
1 0 491 0 0 0 0 312 0 0 0 2
13 25
13 731
2 0 540 0 0 4224 0 324 0 0 981 4
170 303
170 237
190 237
190 232
2 0 569 0 0 0 0 293 0 0 954 3
865 126
869 126
869 169
0 2 569 0 0 0 0 0 316 0 0 4
843 169
1020 169
1020 289
1028 289
4 1 277 0 0 0 0 316 326 0 0 6
1076 271
1149 271
1149 557
716 557
716 339
837 339
4 2 459 0 0 0 0 315 326 0 0 6
1077 317
1134 317
1134 542
730 542
730 348
837 348
4 3 460 0 0 0 0 314 326 0 0 6
1079 360
1119 360
1119 527
745 527
745 357
837 357
4 4 461 0 0 0 0 313 326 0 0 6
1081 404
1107 404
1107 511
758 511
758 366
837 366
1 10 583 0 0 4224 0 316 326 0 0 4
1028 271
919 271
919 366
901 366
1 11 584 0 0 4224 0 315 326 0 0 4
1029 317
914 317
914 375
901 375
1 12 585 0 0 4224 0 314 326 0 0 4
1031 360
909 360
909 384
901 384
13 1 586 0 0 4224 0 326 313 0 0 4
901 393
1025 393
1025 404
1033 404
2 0 569 0 0 0 0 314 0 0 954 3
1031 378
981 378
981 169
2 0 569 0 0 0 0 315 0 0 954 3
1029 335
992 335
992 169
0 2 569 0 0 0 0 0 313 954 0 3
968 169
968 422
1033 422
2 1 587 0 0 8320 0 317 293 0 0 6
833 169
839 169
839 143
827 143
827 126
835 126
1 0 561 0 0 0 0 317 0 0 0 3
803 169
803 168
790 168
3 8 588 0 0 8320 0 324 326 0 0 3
179 348
179 402
837 402
3 7 589 0 0 8320 0 323 326 0 0 3
241 357
241 393
837 393
3 6 590 0 0 8320 0 321 326 0 0 3
313 355
313 384
837 384
3 5 591 0 0 8320 0 319 326 0 0 3
387 355
387 375
837 375
1 0 542 0 0 4096 0 318 0 0 973 3
407 260
407 239
391 239
3 2 542 0 0 4224 0 0 319 0 0 4
391 209
391 302
378 302
378 310
2 1 592 0 0 8320 0 318 319 0 0 4
407 296
407 302
396 302
396 310
1 0 544 0 0 4096 0 320 0 0 976 3
333 260
333 239
317 239
0 2 544 0 0 8320 0 0 321 0 0 5
316 187
317 187
317 302
304 302
304 310
2 1 593 0 0 8320 0 320 321 0 0 4
333 296
333 302
322 302
322 310
1 0 543 0 0 0 0 322 0 0 979 3
261 262
261 241
245 241
3 2 543 0 0 4224 0 0 323 0 0 4
245 211
245 304
232 304
232 312
2 1 594 0 0 8320 0 322 323 0 0 4
261 298
261 304
250 304
250 312
1 0 540 0 0 0 0 325 0 0 0 3
199 253
199 232
183 232
2 1 595 0 0 8320 0 325 324 0 0 4
199 289
199 295
188 295
188 303
16
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
2089 244 2242 292
2102 253 2228 285
7 Digit 1
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 7
758 1674 911 1722
771 1683 897 1715
7 DS-7SEG
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
1060 1581 1269 1629
1074 1589 1254 1621
10 Digit Sort
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 13
1370 1417 1627 1465
1381 1426 1615 1458
13 8-128 Decoder
-16 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 1
384 1760 429 1788
401 1771 411 1791
1 a
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 10
41 536 248 584
54 545 234 577
10 Pull Downs
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 18
721 1249 1068 1297
732 1258 1056 1290
18 Compliment Control
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
1427 853 1846 901
1438 862 1834 894
22 2's compliment creator
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
1552 280 1827 328
1563 289 1815 321
14 System Checker
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 22
920 794 1339 842
931 803 1327 835
22 Bits 4-7 + carry Adder
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
831 429 1108 477
843 437 1095 469
14 Bits 0-3 Adder
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 15
1280 28 1573 76
1291 37 1561 69
15 Toll Programmer
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 8
599 106 766 154
610 115 754 147
8 Displays
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
418 454 693 502
429 463 681 495
14 Pulse Limiters
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 14
175 200 450 248
186 209 438 241
14 Pulse Limiters
-29 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 9
-10 286 175 334
1 294 163 326
9 Selectors
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
